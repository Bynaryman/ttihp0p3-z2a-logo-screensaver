module tt_um_zerotoasic_logo_screensaver (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire \color_index[0] ;
 wire \color_index[1] ;
 wire \color_index[2] ;
 wire dir_x;
 wire dir_y;
 wire \gamepad.decoder.data_reg[0] ;
 wire \gamepad.decoder.data_reg[10] ;
 wire \gamepad.decoder.data_reg[11] ;
 wire \gamepad.decoder.data_reg[1] ;
 wire \gamepad.decoder.data_reg[2] ;
 wire \gamepad.decoder.data_reg[3] ;
 wire \gamepad.decoder.data_reg[4] ;
 wire \gamepad.decoder.data_reg[5] ;
 wire \gamepad.decoder.data_reg[6] ;
 wire \gamepad.decoder.data_reg[7] ;
 wire \gamepad.decoder.data_reg[8] ;
 wire \gamepad.decoder.data_reg[9] ;
 wire \gamepad.driver.pmod_clk_prev ;
 wire \gamepad.driver.pmod_clk_sync[0] ;
 wire \gamepad.driver.pmod_clk_sync[1] ;
 wire \gamepad.driver.pmod_data_sync[0] ;
 wire \gamepad.driver.pmod_data_sync[1] ;
 wire \gamepad.driver.pmod_latch_prev ;
 wire \gamepad.driver.pmod_latch_sync[0] ;
 wire \gamepad.driver.pmod_latch_sync[1] ;
 wire \gamepad.driver.shift_reg[0] ;
 wire \gamepad.driver.shift_reg[10] ;
 wire \gamepad.driver.shift_reg[11] ;
 wire \gamepad.driver.shift_reg[1] ;
 wire \gamepad.driver.shift_reg[2] ;
 wire \gamepad.driver.shift_reg[3] ;
 wire \gamepad.driver.shift_reg[4] ;
 wire \gamepad.driver.shift_reg[5] ;
 wire \gamepad.driver.shift_reg[6] ;
 wire \gamepad.driver.shift_reg[7] ;
 wire \gamepad.driver.shift_reg[8] ;
 wire \gamepad.driver.shift_reg[9] ;
 wire gamepad_start_prev;
 wire hsync;
 wire \logo_left[0] ;
 wire \logo_left[1] ;
 wire \logo_left[2] ;
 wire \logo_left[3] ;
 wire \logo_left[4] ;
 wire \logo_left[5] ;
 wire \logo_left[6] ;
 wire \logo_left[7] ;
 wire \logo_left[8] ;
 wire \logo_left[9] ;
 wire \logo_top[0] ;
 wire \logo_top[1] ;
 wire \logo_top[2] ;
 wire \logo_top[3] ;
 wire \logo_top[4] ;
 wire \logo_top[5] ;
 wire \logo_top[6] ;
 wire \logo_top[7] ;
 wire \logo_top[8] ;
 wire \logo_top[9] ;
 wire manual_mode;
 wire \palette_inst.rrggbb[0] ;
 wire \palette_inst.rrggbb[1] ;
 wire \palette_inst.rrggbb[2] ;
 wire \palette_inst.rrggbb[3] ;
 wire \palette_inst.rrggbb[4] ;
 wire \palette_inst.rrggbb[5] ;
 wire \pix_x[0] ;
 wire \pix_x[1] ;
 wire \pix_x[2] ;
 wire \pix_x[3] ;
 wire \pix_x[4] ;
 wire \pix_x[5] ;
 wire \pix_x[6] ;
 wire \pix_x[7] ;
 wire \pix_x[8] ;
 wire \pix_x[9] ;
 wire \pix_y[0] ;
 wire \pix_y[1] ;
 wire \pix_y[2] ;
 wire \pix_y[3] ;
 wire \pix_y[4] ;
 wire \pix_y[5] ;
 wire \pix_y[6] ;
 wire \pix_y[7] ;
 wire \pix_y[8] ;
 wire \pix_y[9] ;
 wire \prev_y[0] ;
 wire \prev_y[1] ;
 wire \prev_y[2] ;
 wire \prev_y[3] ;
 wire \prev_y[4] ;
 wire \prev_y[5] ;
 wire \prev_y[6] ;
 wire \prev_y[7] ;
 wire \prev_y[8] ;
 wire \prev_y[9] ;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire clknet_0_clk;
 wire \vga_sync_gen.vsync ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;

 sky130_fd_sc_hd__inv_2 _1302_ (.A(\color_index[0] ),
    .Y(_0515_));
 sky130_fd_sc_hd__inv_2 _1303_ (.A(net122),
    .Y(_0516_));
 sky130_fd_sc_hd__inv_2 _1304_ (.A(net124),
    .Y(_0517_));
 sky130_fd_sc_hd__inv_2 _1305_ (.A(dir_x),
    .Y(_0518_));
 sky130_fd_sc_hd__inv_2 _1306_ (.A(\logo_top[8] ),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_2 _1307_ (.A(net125),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _1308_ (.A(net126),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _1309_ (.A(net127),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _1310_ (.A(\logo_left[6] ),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_2 _1311_ (.A(\logo_left[2] ),
    .Y(_0524_));
 sky130_fd_sc_hd__inv_2 _1312_ (.A(net208),
    .Y(_0525_));
 sky130_fd_sc_hd__inv_2 _1313_ (.A(\pix_y[0] ),
    .Y(_0526_));
 sky130_fd_sc_hd__inv_2 _1314_ (.A(net119),
    .Y(_0527_));
 sky130_fd_sc_hd__inv_2 _1315_ (.A(\pix_y[2] ),
    .Y(_0528_));
 sky130_fd_sc_hd__inv_2 _1316_ (.A(\pix_y[3] ),
    .Y(_0529_));
 sky130_fd_sc_hd__inv_2 _1317_ (.A(\pix_y[4] ),
    .Y(_0530_));
 sky130_fd_sc_hd__inv_2 _1318_ (.A(\pix_y[5] ),
    .Y(_0531_));
 sky130_fd_sc_hd__inv_2 _1319_ (.A(net133),
    .Y(_0532_));
 sky130_fd_sc_hd__inv_2 _1320_ (.A(\pix_y[7] ),
    .Y(_0533_));
 sky130_fd_sc_hd__inv_2 _1321_ (.A(\prev_y[1] ),
    .Y(_0534_));
 sky130_fd_sc_hd__inv_2 _1322_ (.A(net3),
    .Y(_0535_));
 sky130_fd_sc_hd__and3_1 _1323_ (.A(\pix_y[5] ),
    .B(\pix_y[6] ),
    .C(\pix_y[7] ),
    .X(_0536_));
 sky130_fd_sc_hd__and4bb_1 _1324_ (.A_N(\pix_y[4] ),
    .B_N(\pix_y[9] ),
    .C(\pix_y[8] ),
    .D(\pix_y[3] ),
    .X(_0537_));
 sky130_fd_sc_hd__and4_1 _1325_ (.A(\pix_y[1] ),
    .B(_0528_),
    .C(_0536_),
    .D(_0537_),
    .X(_0005_));
 sky130_fd_sc_hd__or3_1 _1326_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(\pix_x[6] ),
    .X(_0538_));
 sky130_fd_sc_hd__a31oi_1 _1327_ (.A1(\pix_x[4] ),
    .A2(\pix_x[5] ),
    .A3(\pix_x[6] ),
    .B1(\pix_x[8] ),
    .Y(_0539_));
 sky130_fd_sc_hd__and4_1 _1328_ (.A(\pix_x[7] ),
    .B(\pix_x[9] ),
    .C(_0538_),
    .D(_0539_),
    .X(_0004_));
 sky130_fd_sc_hd__xnor2_1 _1329_ (.A(\pix_y[9] ),
    .B(\prev_y[9] ),
    .Y(_0540_));
 sky130_fd_sc_hd__xnor2_1 _1330_ (.A(net118),
    .B(\prev_y[8] ),
    .Y(_0541_));
 sky130_fd_sc_hd__xor2_1 _1331_ (.A(\pix_y[5] ),
    .B(\prev_y[5] ),
    .X(_0542_));
 sky130_fd_sc_hd__a221oi_1 _1332_ (.A1(_0528_),
    .A2(\prev_y[2] ),
    .B1(\prev_y[3] ),
    .B2(_0529_),
    .C1(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__xnor2_1 _1333_ (.A(\pix_y[6] ),
    .B(\prev_y[6] ),
    .Y(_0544_));
 sky130_fd_sc_hd__o2bb2a_1 _1334_ (.A1_N(_0530_),
    .A2_N(\prev_y[4] ),
    .B1(\prev_y[3] ),
    .B2(_0529_),
    .X(_0545_));
 sky130_fd_sc_hd__o221a_1 _1335_ (.A1(_0527_),
    .A2(\prev_y[1] ),
    .B1(\prev_y[7] ),
    .B2(_0533_),
    .C1(_0541_),
    .X(_0546_));
 sky130_fd_sc_hd__a22oi_1 _1336_ (.A1(_0526_),
    .A2(\prev_y[0] ),
    .B1(\prev_y[7] ),
    .B2(_0533_),
    .Y(_0547_));
 sky130_fd_sc_hd__o221a_1 _1337_ (.A1(_0526_),
    .A2(\prev_y[0] ),
    .B1(_0534_),
    .B2(net119),
    .C1(_0545_),
    .X(_0548_));
 sky130_fd_sc_hd__o221a_1 _1338_ (.A1(_0528_),
    .A2(\prev_y[2] ),
    .B1(\prev_y[4] ),
    .B2(_0530_),
    .C1(_0547_),
    .X(_0549_));
 sky130_fd_sc_hd__and4_1 _1339_ (.A(_0540_),
    .B(_0544_),
    .C(_0548_),
    .D(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__or4_1 _1340_ (.A(\pix_y[4] ),
    .B(\pix_y[5] ),
    .C(\pix_y[6] ),
    .D(\pix_y[7] ),
    .X(_0551_));
 sky130_fd_sc_hd__or4_1 _1341_ (.A(\pix_y[0] ),
    .B(net119),
    .C(\pix_y[2] ),
    .D(\pix_y[9] ),
    .X(_0552_));
 sky130_fd_sc_hd__or4_1 _1342_ (.A(\pix_y[3] ),
    .B(net118),
    .C(_0551_),
    .D(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__a31o_4 _1343_ (.A1(_0543_),
    .A2(_0546_),
    .A3(_0550_),
    .B1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__or2_1 _1344_ (.A(net120),
    .B(_0554_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _1345_ (.A(\logo_top[1] ),
    .B(\logo_top[0] ),
    .Y(_0556_));
 sky130_fd_sc_hd__and3_1 _1346_ (.A(\logo_top[2] ),
    .B(\logo_top[1] ),
    .C(\logo_top[0] ),
    .X(_0557_));
 sky130_fd_sc_hd__and3_1 _1347_ (.A(net128),
    .B(net129),
    .C(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__and4_1 _1348_ (.A(net125),
    .B(net126),
    .C(\logo_top[5] ),
    .D(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__xnor2_1 _1349_ (.A(_0519_),
    .B(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__or2_1 _1350_ (.A(\logo_top[9] ),
    .B(net125),
    .X(_0561_));
 sky130_fd_sc_hd__nor2_1 _1351_ (.A(_0521_),
    .B(_0561_),
    .Y(_0562_));
 sky130_fd_sc_hd__and4_1 _1352_ (.A(\logo_top[8] ),
    .B(_0522_),
    .C(_0558_),
    .D(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__nand2_1 _1353_ (.A(dir_y),
    .B(_0563_),
    .Y(_0564_));
 sky130_fd_sc_hd__or2_1 _1354_ (.A(net129),
    .B(\logo_top[2] ),
    .X(_0565_));
 sky130_fd_sc_hd__nor2_1 _1355_ (.A(net127),
    .B(net128),
    .Y(_0566_));
 sky130_fd_sc_hd__or3_1 _1356_ (.A(net127),
    .B(net128),
    .C(_0565_),
    .X(_0567_));
 sky130_fd_sc_hd__nor2_1 _1357_ (.A(net126),
    .B(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__or2_1 _1358_ (.A(dir_y),
    .B(\logo_top[8] ),
    .X(_0569_));
 sky130_fd_sc_hd__or2_1 _1359_ (.A(\logo_left[5] ),
    .B(net130),
    .X(_0570_));
 sky130_fd_sc_hd__or3_1 _1360_ (.A(\logo_left[6] ),
    .B(net131),
    .C(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__or3b_1 _1361_ (.A(\logo_left[2] ),
    .B(\logo_left[1] ),
    .C_N(\logo_left[0] ),
    .X(_0572_));
 sky130_fd_sc_hd__or2_1 _1362_ (.A(dir_x),
    .B(\logo_left[9] ),
    .X(_0573_));
 sky130_fd_sc_hd__or2_1 _1363_ (.A(\logo_left[8] ),
    .B(\logo_left[7] ),
    .X(_0574_));
 sky130_fd_sc_hd__or4_1 _1364_ (.A(_0571_),
    .B(_0572_),
    .C(_0573_),
    .D(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nand2_1 _1365_ (.A(\logo_left[1] ),
    .B(\logo_left[0] ),
    .Y(_0576_));
 sky130_fd_sc_hd__nor2_1 _1366_ (.A(_0524_),
    .B(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__and3_1 _1367_ (.A(\logo_left[5] ),
    .B(net130),
    .C(net131),
    .X(_0578_));
 sky130_fd_sc_hd__and4_1 _1368_ (.A(\logo_left[7] ),
    .B(\logo_left[6] ),
    .C(_0577_),
    .D(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__and2_1 _1369_ (.A(\logo_left[8] ),
    .B(_0579_),
    .X(_0580_));
 sky130_fd_sc_hd__or3b_1 _1370_ (.A(net126),
    .B(\logo_top[1] ),
    .C_N(\logo_top[0] ),
    .X(_0581_));
 sky130_fd_sc_hd__or4_1 _1371_ (.A(_0561_),
    .B(_0567_),
    .C(_0569_),
    .D(_0581_),
    .X(_0582_));
 sky130_fd_sc_hd__or4_1 _1372_ (.A(\logo_left[6] ),
    .B(net131),
    .C(_0572_),
    .D(_0574_),
    .X(_0583_));
 sky130_fd_sc_hd__nand2_1 _1373_ (.A(dir_x),
    .B(_0580_),
    .Y(_0584_));
 sky130_fd_sc_hd__o32a_1 _1374_ (.A1(_0570_),
    .A2(_0573_),
    .A3(_0583_),
    .B1(_0584_),
    .B2(\logo_left[9] ),
    .X(_0585_));
 sky130_fd_sc_hd__a31o_1 _1375_ (.A1(_0564_),
    .A2(_0582_),
    .A3(_0585_),
    .B1(_0555_),
    .X(_0586_));
 sky130_fd_sc_hd__or4_1 _1376_ (.A(_0561_),
    .B(_0567_),
    .C(_0569_),
    .D(_0581_),
    .X(_0587_));
 sky130_fd_sc_hd__and2_1 _1377_ (.A(_0515_),
    .B(_0586_),
    .X(_0588_));
 sky130_fd_sc_hd__nor2_1 _1378_ (.A(_0515_),
    .B(_0586_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor2_1 _1379_ (.A(_0588_),
    .B(_0589_),
    .Y(_0590_));
 sky130_fd_sc_hd__nand2_1 _1380_ (.A(net135),
    .B(_0590_),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_2 _1381_ (.A(_0591_),
    .Y(_0054_));
 sky130_fd_sc_hd__nand2_1 _1382_ (.A(\color_index[1] ),
    .B(_0589_),
    .Y(_0592_));
 sky130_fd_sc_hd__xnor2_1 _1383_ (.A(\color_index[2] ),
    .B(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a21o_1 _1384_ (.A1(net206),
    .A2(_0593_),
    .B1(_0591_),
    .X(_0000_));
 sky130_fd_sc_hd__or2_1 _1385_ (.A(\color_index[1] ),
    .B(_0589_),
    .X(_0594_));
 sky130_fd_sc_hd__and3_1 _1386_ (.A(net135),
    .B(_0592_),
    .C(_0594_),
    .X(_0055_));
 sky130_fd_sc_hd__nand2_1 _1387_ (.A(net135),
    .B(_0593_),
    .Y(_0595_));
 sky130_fd_sc_hd__inv_2 _1388_ (.A(_0595_),
    .Y(_0056_));
 sky130_fd_sc_hd__and2_1 _1389_ (.A(_0054_),
    .B(_0593_),
    .X(_0596_));
 sky130_fd_sc_hd__xnor2_1 _1390_ (.A(_0055_),
    .B(_0596_),
    .Y(_0001_));
 sky130_fd_sc_hd__nand2_1 _1391_ (.A(_0591_),
    .B(_0595_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1392_ (.A(_0100_),
    .Y(_0597_));
 sky130_fd_sc_hd__nor3_1 _1393_ (.A(\color_index[2] ),
    .B(\color_index[1] ),
    .C(_0591_),
    .Y(_0598_));
 sky130_fd_sc_hd__a211o_1 _1394_ (.A1(_0055_),
    .A2(_0597_),
    .B1(_0598_),
    .C1(_0596_),
    .X(_0002_));
 sky130_fd_sc_hd__o21ba_1 _1395_ (.A1(_0590_),
    .A2(_0595_),
    .B1_N(_0598_),
    .X(_0003_));
 sky130_fd_sc_hd__nand2b_2 _1396_ (.A_N(\pix_x[0] ),
    .B(\logo_left[0] ),
    .Y(_0599_));
 sky130_fd_sc_hd__and2b_1 _1397_ (.A_N(\logo_left[1] ),
    .B(\pix_x[1] ),
    .X(_0600_));
 sky130_fd_sc_hd__xnor2_2 _1398_ (.A(\logo_left[1] ),
    .B(\pix_x[1] ),
    .Y(_0601_));
 sky130_fd_sc_hd__xor2_2 _1399_ (.A(_0599_),
    .B(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__and2_1 _1400_ (.A(_0521_),
    .B(\pix_y[6] ),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_1 _1401_ (.A(_0521_),
    .B(\pix_y[6] ),
    .Y(_0604_));
 sky130_fd_sc_hd__nor2_2 _1402_ (.A(_0603_),
    .B(_0604_),
    .Y(_0605_));
 sky130_fd_sc_hd__nor2_1 _1403_ (.A(net128),
    .B(_0530_),
    .Y(_0606_));
 sky130_fd_sc_hd__nor2_1 _1404_ (.A(net129),
    .B(_0529_),
    .Y(_0607_));
 sky130_fd_sc_hd__and2_1 _1405_ (.A(net129),
    .B(_0529_),
    .X(_0608_));
 sky130_fd_sc_hd__or2_2 _1406_ (.A(_0607_),
    .B(_0608_),
    .X(_0609_));
 sky130_fd_sc_hd__and2b_1 _1407_ (.A_N(\logo_top[2] ),
    .B(\pix_y[2] ),
    .X(_0610_));
 sky130_fd_sc_hd__and2b_1 _1408_ (.A_N(\logo_top[1] ),
    .B(net119),
    .X(_0611_));
 sky130_fd_sc_hd__nand2b_2 _1409_ (.A_N(\pix_y[0] ),
    .B(\logo_top[0] ),
    .Y(_0612_));
 sky130_fd_sc_hd__xnor2_4 _1410_ (.A(\logo_top[1] ),
    .B(net119),
    .Y(_0613_));
 sky130_fd_sc_hd__a21o_2 _1411_ (.A1(_0612_),
    .A2(_0613_),
    .B1(_0611_),
    .X(_0614_));
 sky130_fd_sc_hd__and2b_1 _1412_ (.A_N(\pix_y[2] ),
    .B(\logo_top[2] ),
    .X(_0615_));
 sky130_fd_sc_hd__nor2_2 _1413_ (.A(_0610_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__a21oi_4 _1414_ (.A1(_0614_),
    .A2(_0616_),
    .B1(_0610_),
    .Y(_0617_));
 sky130_fd_sc_hd__o21bai_4 _1415_ (.A1(_0608_),
    .A2(_0617_),
    .B1_N(_0607_),
    .Y(_0618_));
 sky130_fd_sc_hd__and2_1 _1416_ (.A(\logo_top[4] ),
    .B(_0530_),
    .X(_0619_));
 sky130_fd_sc_hd__nor2_2 _1417_ (.A(_0606_),
    .B(_0619_),
    .Y(_0620_));
 sky130_fd_sc_hd__a21o_1 _1418_ (.A1(_0618_),
    .A2(_0620_),
    .B1(_0606_),
    .X(_0621_));
 sky130_fd_sc_hd__a21oi_1 _1419_ (.A1(_0522_),
    .A2(\pix_y[5] ),
    .B1(_0621_),
    .Y(_0622_));
 sky130_fd_sc_hd__a21oi_4 _1420_ (.A1(net127),
    .A2(_0531_),
    .B1(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__xor2_2 _1421_ (.A(_0605_),
    .B(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__xnor2_4 _1422_ (.A(_0605_),
    .B(_0623_),
    .Y(_0625_));
 sky130_fd_sc_hd__xor2_2 _1423_ (.A(_0609_),
    .B(_0617_),
    .X(_0626_));
 sky130_fd_sc_hd__xnor2_4 _1424_ (.A(_0609_),
    .B(_0617_),
    .Y(_0627_));
 sky130_fd_sc_hd__xor2_1 _1425_ (.A(_0614_),
    .B(_0616_),
    .X(_0628_));
 sky130_fd_sc_hd__xnor2_2 _1426_ (.A(_0614_),
    .B(_0616_),
    .Y(_0629_));
 sky130_fd_sc_hd__nor2_4 _1427_ (.A(net85),
    .B(net99),
    .Y(_0630_));
 sky130_fd_sc_hd__nand2_1 _1428_ (.A(net81),
    .B(net102),
    .Y(_0631_));
 sky130_fd_sc_hd__xor2_2 _1429_ (.A(_0612_),
    .B(_0613_),
    .X(_0632_));
 sky130_fd_sc_hd__xnor2_1 _1430_ (.A(_0612_),
    .B(_0613_),
    .Y(_0633_));
 sky130_fd_sc_hd__and2_1 _1431_ (.A(_0523_),
    .B(\pix_x[6] ),
    .X(_0634_));
 sky130_fd_sc_hd__nor2_1 _1432_ (.A(_0523_),
    .B(\pix_x[6] ),
    .Y(_0635_));
 sky130_fd_sc_hd__nor2_1 _1433_ (.A(_0634_),
    .B(_0635_),
    .Y(_0636_));
 sky130_fd_sc_hd__and2b_1 _1434_ (.A_N(\pix_x[5] ),
    .B(\logo_left[5] ),
    .X(_0637_));
 sky130_fd_sc_hd__nand2b_1 _1435_ (.A_N(\pix_x[5] ),
    .B(\logo_left[5] ),
    .Y(_0638_));
 sky130_fd_sc_hd__and2b_1 _1436_ (.A_N(\logo_left[5] ),
    .B(\pix_x[5] ),
    .X(_0639_));
 sky130_fd_sc_hd__and2b_1 _1437_ (.A_N(net130),
    .B(\pix_x[4] ),
    .X(_0640_));
 sky130_fd_sc_hd__and2b_1 _1438_ (.A_N(\pix_x[4] ),
    .B(net130),
    .X(_0641_));
 sky130_fd_sc_hd__nor2_2 _1439_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__and2b_1 _1440_ (.A_N(\logo_left[2] ),
    .B(\pix_x[2] ),
    .X(_0643_));
 sky130_fd_sc_hd__and2b_1 _1441_ (.A_N(\pix_x[2] ),
    .B(\logo_left[2] ),
    .X(_0644_));
 sky130_fd_sc_hd__nor2_2 _1442_ (.A(_0643_),
    .B(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__a21o_2 _1443_ (.A1(_0599_),
    .A2(_0601_),
    .B1(_0600_),
    .X(_0646_));
 sky130_fd_sc_hd__and2b_1 _1444_ (.A_N(net131),
    .B(\pix_x[3] ),
    .X(_0647_));
 sky130_fd_sc_hd__xnor2_4 _1445_ (.A(net131),
    .B(\pix_x[3] ),
    .Y(_0648_));
 sky130_fd_sc_hd__a31o_1 _1446_ (.A1(_0524_),
    .A2(\pix_x[2] ),
    .A3(_0648_),
    .B1(_0647_),
    .X(_0649_));
 sky130_fd_sc_hd__a31o_2 _1447_ (.A1(_0645_),
    .A2(_0646_),
    .A3(_0648_),
    .B1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__a21o_1 _1448_ (.A1(_0642_),
    .A2(_0650_),
    .B1(_0640_),
    .X(_0651_));
 sky130_fd_sc_hd__a211o_1 _1449_ (.A1(_0642_),
    .A2(_0650_),
    .B1(_0639_),
    .C1(_0640_),
    .X(_0652_));
 sky130_fd_sc_hd__and3_1 _1450_ (.A(_0636_),
    .B(_0638_),
    .C(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nand3_2 _1451_ (.A(_0636_),
    .B(_0638_),
    .C(_0652_),
    .Y(_0654_));
 sky130_fd_sc_hd__a21oi_2 _1452_ (.A1(_0638_),
    .A2(_0652_),
    .B1(_0636_),
    .Y(_0655_));
 sky130_fd_sc_hd__a21o_2 _1453_ (.A1(_0638_),
    .A2(_0652_),
    .B1(_0636_),
    .X(_0656_));
 sky130_fd_sc_hd__nor2_1 _1454_ (.A(net65),
    .B(net59),
    .Y(_0657_));
 sky130_fd_sc_hd__nand2_1 _1455_ (.A(net60),
    .B(net55),
    .Y(_0658_));
 sky130_fd_sc_hd__nor2_1 _1456_ (.A(_0637_),
    .B(_0639_),
    .Y(_0659_));
 sky130_fd_sc_hd__xnor2_1 _1457_ (.A(_0651_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__xor2_1 _1458_ (.A(_0651_),
    .B(_0659_),
    .X(_0661_));
 sky130_fd_sc_hd__and3_2 _1459_ (.A(net60),
    .B(net55),
    .C(net45),
    .X(_0662_));
 sky130_fd_sc_hd__or3_1 _1460_ (.A(net64),
    .B(net58),
    .C(net52),
    .X(_0663_));
 sky130_fd_sc_hd__xor2_2 _1461_ (.A(_0642_),
    .B(_0650_),
    .X(_0664_));
 sky130_fd_sc_hd__xnor2_1 _1462_ (.A(_0642_),
    .B(_0650_),
    .Y(_0665_));
 sky130_fd_sc_hd__nand2_1 _1463_ (.A(net46),
    .B(net77),
    .Y(_0666_));
 sky130_fd_sc_hd__o22a_1 _1464_ (.A1(net63),
    .A2(net59),
    .B1(net53),
    .B2(net79),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_2 _1465_ (.A1(net61),
    .A2(net56),
    .B1(net48),
    .B2(net78),
    .X(_0668_));
 sky130_fd_sc_hd__nor2_1 _1466_ (.A(net23),
    .B(net44),
    .Y(_0669_));
 sky130_fd_sc_hd__or3_4 _1467_ (.A(net64),
    .B(net58),
    .C(net44),
    .X(_0670_));
 sky130_fd_sc_hd__o211a_1 _1468_ (.A1(net63),
    .A2(net59),
    .B1(net47),
    .C1(net77),
    .X(_0671_));
 sky130_fd_sc_hd__a211o_1 _1469_ (.A1(net61),
    .A2(net57),
    .B1(net53),
    .C1(net79),
    .X(_0672_));
 sky130_fd_sc_hd__nor2_1 _1470_ (.A(_0662_),
    .B(net21),
    .Y(_0673_));
 sky130_fd_sc_hd__a21oi_4 _1471_ (.A1(_0645_),
    .A2(_0646_),
    .B1(_0643_),
    .Y(_0674_));
 sky130_fd_sc_hd__xor2_4 _1472_ (.A(_0648_),
    .B(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__xnor2_2 _1473_ (.A(_0648_),
    .B(_0674_),
    .Y(_0676_));
 sky130_fd_sc_hd__nor2_1 _1474_ (.A(net50),
    .B(net76),
    .Y(_0677_));
 sky130_fd_sc_hd__nand2_1 _1475_ (.A(net48),
    .B(net75),
    .Y(_0678_));
 sky130_fd_sc_hd__nor2_1 _1476_ (.A(net28),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__a211o_2 _1477_ (.A1(net60),
    .A2(net55),
    .B1(net51),
    .C1(net76),
    .X(_0680_));
 sky130_fd_sc_hd__o211a_1 _1478_ (.A1(_0662_),
    .A2(net21),
    .B1(_0680_),
    .C1(net111),
    .X(_0681_));
 sky130_fd_sc_hd__nand2_1 _1479_ (.A(net47),
    .B(net79),
    .Y(_0682_));
 sky130_fd_sc_hd__or2_1 _1480_ (.A(\logo_top[0] ),
    .B(_0526_),
    .X(_0683_));
 sky130_fd_sc_hd__and2_2 _1481_ (.A(_0612_),
    .B(_0683_),
    .X(_0684_));
 sky130_fd_sc_hd__nand2_2 _1482_ (.A(_0612_),
    .B(_0683_),
    .Y(_0685_));
 sky130_fd_sc_hd__nor2_1 _1483_ (.A(net112),
    .B(net90),
    .Y(_0686_));
 sky130_fd_sc_hd__nand2_2 _1484_ (.A(_0613_),
    .B(net94),
    .Y(_0687_));
 sky130_fd_sc_hd__nor2_1 _1485_ (.A(net78),
    .B(net76),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_4 _1486_ (.A(net80),
    .B(net75),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _1487_ (.A(net51),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__o22a_2 _1488_ (.A1(net64),
    .A2(net58),
    .B1(net46),
    .B2(net43),
    .X(_0691_));
 sky130_fd_sc_hd__a22o_1 _1489_ (.A1(net62),
    .A2(net57),
    .B1(net50),
    .B2(_0689_),
    .X(_0692_));
 sky130_fd_sc_hd__a21o_2 _1490_ (.A1(net62),
    .A2(net56),
    .B1(net46),
    .X(_0693_));
 sky130_fd_sc_hd__a211o_2 _1491_ (.A1(net60),
    .A2(net55),
    .B1(net45),
    .C1(net43),
    .X(_0694_));
 sky130_fd_sc_hd__nand2_1 _1492_ (.A(_0670_),
    .B(_0692_),
    .Y(_0695_));
 sky130_fd_sc_hd__a31oi_1 _1493_ (.A1(net22),
    .A2(net20),
    .A3(_0694_),
    .B1(net73),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_1 _1494_ (.A(net112),
    .B(net94),
    .Y(_0697_));
 sky130_fd_sc_hd__or2_4 _1495_ (.A(net112),
    .B(net94),
    .X(_0698_));
 sky130_fd_sc_hd__nor2_4 _1496_ (.A(net77),
    .B(net75),
    .Y(_0699_));
 sky130_fd_sc_hd__o22a_2 _1497_ (.A1(net63),
    .A2(net59),
    .B1(net44),
    .B2(net79),
    .X(_0700_));
 sky130_fd_sc_hd__a221o_1 _1498_ (.A1(_0654_),
    .A2(_0656_),
    .B1(net51),
    .B2(net78),
    .C1(_0699_),
    .X(_0701_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(_0670_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__and3_1 _1500_ (.A(_0670_),
    .B(_0697_),
    .C(_0701_),
    .X(_0703_));
 sky130_fd_sc_hd__o31a_1 _1501_ (.A1(_0681_),
    .A2(_0696_),
    .A3(_0703_),
    .B1(_0630_),
    .X(_0704_));
 sky130_fd_sc_hd__xor2_4 _1502_ (.A(_0618_),
    .B(_0620_),
    .X(_0705_));
 sky130_fd_sc_hd__xnor2_1 _1503_ (.A(_0618_),
    .B(_0620_),
    .Y(_0706_));
 sky130_fd_sc_hd__nor2_1 _1504_ (.A(net46),
    .B(_0689_),
    .Y(_0707_));
 sky130_fd_sc_hd__nor2_8 _1505_ (.A(net80),
    .B(net75),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_4 _1506_ (.A(net77),
    .B(_0675_),
    .Y(_0709_));
 sky130_fd_sc_hd__nor2_2 _1507_ (.A(net51),
    .B(_0708_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_4 _1508_ (.A(net48),
    .B(_0709_),
    .Y(_0711_));
 sky130_fd_sc_hd__or4_1 _1509_ (.A(net64),
    .B(net58),
    .C(net52),
    .D(_0708_),
    .X(_0712_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(_0668_),
    .B(_0712_),
    .Y(_0713_));
 sky130_fd_sc_hd__xnor2_4 _1511_ (.A(net54),
    .B(net79),
    .Y(_0714_));
 sky130_fd_sc_hd__inv_2 _1512_ (.A(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__mux2_1 _1513_ (.A0(net77),
    .A1(net43),
    .S(net52),
    .X(_0716_));
 sky130_fd_sc_hd__o21ai_2 _1514_ (.A1(net28),
    .A2(_0716_),
    .B1(net18),
    .Y(_0717_));
 sky130_fd_sc_hd__o21a_1 _1515_ (.A1(net28),
    .A2(_0716_),
    .B1(net18),
    .X(_0718_));
 sky130_fd_sc_hd__nor2_1 _1516_ (.A(net86),
    .B(net100),
    .Y(_0719_));
 sky130_fd_sc_hd__nand2_2 _1517_ (.A(net81),
    .B(net98),
    .Y(_0720_));
 sky130_fd_sc_hd__a21oi_1 _1518_ (.A1(_0717_),
    .A2(net35),
    .B1(net38),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_2 _1519_ (.A(net46),
    .B(net43),
    .Y(_0722_));
 sky130_fd_sc_hd__inv_2 _1520_ (.A(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__o211a_1 _1521_ (.A1(net64),
    .A2(net58),
    .B1(net45),
    .C1(net43),
    .X(_0724_));
 sky130_fd_sc_hd__a211o_2 _1522_ (.A1(net62),
    .A2(net57),
    .B1(net52),
    .C1(_0689_),
    .X(_0725_));
 sky130_fd_sc_hd__and3_1 _1523_ (.A(net60),
    .B(net55),
    .C(net78),
    .X(_0726_));
 sky130_fd_sc_hd__or3_4 _1524_ (.A(net63),
    .B(net59),
    .C(net79),
    .X(_0727_));
 sky130_fd_sc_hd__and4_2 _1525_ (.A(net60),
    .B(net55),
    .C(net50),
    .D(net78),
    .X(_0728_));
 sky130_fd_sc_hd__or2_1 _1526_ (.A(_0724_),
    .B(_0728_),
    .X(_0729_));
 sky130_fd_sc_hd__nor2_1 _1527_ (.A(net108),
    .B(net94),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_1 _1528_ (.A(net105),
    .B(net94),
    .X(_0731_));
 sky130_fd_sc_hd__o211a_4 _1529_ (.A1(net48),
    .A2(_0709_),
    .B1(net62),
    .C1(net57),
    .X(_0732_));
 sky130_fd_sc_hd__a211o_1 _1530_ (.A1(net50),
    .A2(_0708_),
    .B1(net64),
    .C1(net58),
    .X(_0733_));
 sky130_fd_sc_hd__a22o_1 _1531_ (.A1(net60),
    .A2(net55),
    .B1(net44),
    .B2(_0688_),
    .X(_0734_));
 sky130_fd_sc_hd__nand2_1 _1532_ (.A(_0733_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__a21o_1 _1533_ (.A1(_0733_),
    .A2(_0734_),
    .B1(net69),
    .X(_0736_));
 sky130_fd_sc_hd__nor2_1 _1534_ (.A(net83),
    .B(net99),
    .Y(_0737_));
 sky130_fd_sc_hd__nand2_1 _1535_ (.A(net85),
    .B(net100),
    .Y(_0738_));
 sky130_fd_sc_hd__a21oi_1 _1536_ (.A1(_0729_),
    .A2(_0736_),
    .B1(net32),
    .Y(_0739_));
 sky130_fd_sc_hd__nor2_4 _1537_ (.A(net81),
    .B(net100),
    .Y(_0740_));
 sky130_fd_sc_hd__nand2_2 _1538_ (.A(net86),
    .B(net99),
    .Y(_0741_));
 sky130_fd_sc_hd__and3_2 _1539_ (.A(net61),
    .B(net56),
    .C(_0689_),
    .X(_0742_));
 sky130_fd_sc_hd__or2_1 _1540_ (.A(net24),
    .B(_0690_),
    .X(_0743_));
 sky130_fd_sc_hd__o21ai_1 _1541_ (.A1(net24),
    .A2(_0690_),
    .B1(_0725_),
    .Y(_0744_));
 sky130_fd_sc_hd__o211a_1 _1542_ (.A1(net24),
    .A2(_0690_),
    .B1(_0725_),
    .C1(net111),
    .X(_0745_));
 sky130_fd_sc_hd__inv_2 _1543_ (.A(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__and3_2 _1544_ (.A(net60),
    .B(net55),
    .C(net43),
    .X(_0747_));
 sky130_fd_sc_hd__or3_2 _1545_ (.A(net64),
    .B(net58),
    .C(_0689_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _1546_ (.A(net97),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__nand2_1 _1547_ (.A(net77),
    .B(net75),
    .Y(_0750_));
 sky130_fd_sc_hd__xnor2_4 _1548_ (.A(net78),
    .B(net76),
    .Y(_0751_));
 sky130_fd_sc_hd__xnor2_4 _1549_ (.A(net79),
    .B(_0675_),
    .Y(_0752_));
 sky130_fd_sc_hd__nand2_1 _1550_ (.A(net44),
    .B(_0751_),
    .Y(_0753_));
 sky130_fd_sc_hd__a21o_2 _1551_ (.A1(net61),
    .A2(net56),
    .B1(_0752_),
    .X(_0754_));
 sky130_fd_sc_hd__o21a_1 _1552_ (.A1(net51),
    .A2(_0754_),
    .B1(_0670_),
    .X(_0755_));
 sky130_fd_sc_hd__o31a_1 _1553_ (.A1(_0745_),
    .A2(_0749_),
    .A3(_0755_),
    .B1(_0740_),
    .X(_0756_));
 sky130_fd_sc_hd__or4b_1 _1554_ (.A(_0704_),
    .B(_0739_),
    .C(_0756_),
    .D_N(_0721_),
    .X(_0757_));
 sky130_fd_sc_hd__xnor2_1 _1555_ (.A(net127),
    .B(\pix_y[5] ),
    .Y(_0758_));
 sky130_fd_sc_hd__xnor2_1 _1556_ (.A(_0621_),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__xor2_1 _1557_ (.A(_0621_),
    .B(_0758_),
    .X(_0760_));
 sky130_fd_sc_hd__nor2_4 _1558_ (.A(net48),
    .B(_0708_),
    .Y(_0761_));
 sky130_fd_sc_hd__nand2_4 _1559_ (.A(net52),
    .B(_0709_),
    .Y(_0762_));
 sky130_fd_sc_hd__nand2_1 _1560_ (.A(net47),
    .B(_0752_),
    .Y(_0763_));
 sky130_fd_sc_hd__and3_1 _1561_ (.A(net74),
    .B(_0753_),
    .C(_0762_),
    .X(_0764_));
 sky130_fd_sc_hd__o211a_1 _1562_ (.A1(net64),
    .A2(net58),
    .B1(net50),
    .C1(net78),
    .X(_0765_));
 sky130_fd_sc_hd__a211o_1 _1563_ (.A1(net62),
    .A2(net57),
    .B1(net48),
    .C1(net80),
    .X(_0766_));
 sky130_fd_sc_hd__and2_2 _1564_ (.A(net18),
    .B(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__and3_1 _1565_ (.A(net18),
    .B(_0725_),
    .C(_0766_),
    .X(_0768_));
 sky130_fd_sc_hd__nand2_1 _1566_ (.A(net47),
    .B(net76),
    .Y(_0769_));
 sky130_fd_sc_hd__o22a_1 _1567_ (.A1(net65),
    .A2(_0655_),
    .B1(net52),
    .B2(net77),
    .X(_0770_));
 sky130_fd_sc_hd__xnor2_2 _1568_ (.A(net50),
    .B(net76),
    .Y(_0771_));
 sky130_fd_sc_hd__xnor2_2 _1569_ (.A(net44),
    .B(net76),
    .Y(_0772_));
 sky130_fd_sc_hd__or3_1 _1570_ (.A(net28),
    .B(net80),
    .C(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__nor2_1 _1571_ (.A(net69),
    .B(_0768_),
    .Y(_0774_));
 sky130_fd_sc_hd__a21oi_1 _1572_ (.A1(net18),
    .A2(_0773_),
    .B1(net71),
    .Y(_0775_));
 sky130_fd_sc_hd__o31a_1 _1573_ (.A1(_0764_),
    .A2(_0774_),
    .A3(_0775_),
    .B1(_0630_),
    .X(_0776_));
 sky130_fd_sc_hd__nor2_4 _1574_ (.A(net101),
    .B(net111),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2_4 _1575_ (.A(net99),
    .B(net107),
    .Y(_0778_));
 sky130_fd_sc_hd__o21a_2 _1576_ (.A1(net28),
    .A2(_0714_),
    .B1(net18),
    .X(_0779_));
 sky130_fd_sc_hd__o21ai_1 _1577_ (.A1(_0777_),
    .A2(_0779_),
    .B1(_0768_),
    .Y(_0780_));
 sky130_fd_sc_hd__a21oi_1 _1578_ (.A1(net87),
    .A2(_0780_),
    .B1(net42),
    .Y(_0781_));
 sky130_fd_sc_hd__a21o_1 _1579_ (.A1(net87),
    .A2(_0780_),
    .B1(net42),
    .X(_0782_));
 sky130_fd_sc_hd__or2_1 _1580_ (.A(net45),
    .B(net30),
    .X(_0783_));
 sky130_fd_sc_hd__o22a_1 _1581_ (.A1(net63),
    .A2(net59),
    .B1(net46),
    .B2(net30),
    .X(_0784_));
 sky130_fd_sc_hd__a2bb2o_2 _1582_ (.A1_N(net44),
    .A2_N(net30),
    .B1(net61),
    .B2(net56),
    .X(_0785_));
 sky130_fd_sc_hd__a21oi_4 _1583_ (.A1(net53),
    .A2(net75),
    .B1(_0699_),
    .Y(_0786_));
 sky130_fd_sc_hd__a21oi_1 _1584_ (.A1(net26),
    .A2(_0786_),
    .B1(_0784_),
    .Y(_0787_));
 sky130_fd_sc_hd__a21o_1 _1585_ (.A1(net26),
    .A2(_0786_),
    .B1(_0784_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _1586_ (.A(net44),
    .B(_0708_),
    .Y(_0789_));
 sky130_fd_sc_hd__xnor2_4 _1587_ (.A(net52),
    .B(_0708_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_1 _1588_ (.A(net24),
    .B(_0790_),
    .Y(_0791_));
 sky130_fd_sc_hd__o2bb2a_1 _1589_ (.A1_N(net24),
    .A2_N(_0790_),
    .B1(_0699_),
    .B2(net22),
    .X(_0792_));
 sky130_fd_sc_hd__a2bb2o_1 _1590_ (.A1_N(_0792_),
    .A2_N(_0698_),
    .B1(net74),
    .B2(_0788_),
    .X(_0793_));
 sky130_fd_sc_hd__a21o_1 _1591_ (.A1(net53),
    .A2(_0689_),
    .B1(_0752_),
    .X(_0794_));
 sky130_fd_sc_hd__nand2_1 _1592_ (.A(_0691_),
    .B(_0751_),
    .Y(_0795_));
 sky130_fd_sc_hd__and3_1 _1593_ (.A(net71),
    .B(_0762_),
    .C(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__nor2_4 _1594_ (.A(net108),
    .B(net91),
    .Y(_0797_));
 sky130_fd_sc_hd__nand2_8 _1595_ (.A(net112),
    .B(net94),
    .Y(_0798_));
 sky130_fd_sc_hd__nor2_1 _1596_ (.A(_0792_),
    .B(_0798_),
    .Y(_0799_));
 sky130_fd_sc_hd__o31a_1 _1597_ (.A1(_0793_),
    .A2(_0796_),
    .A3(_0799_),
    .B1(net35),
    .X(_0800_));
 sky130_fd_sc_hd__o311a_1 _1598_ (.A1(_0776_),
    .A2(_0782_),
    .A3(_0800_),
    .B1(net13),
    .C1(_0757_),
    .X(_0801_));
 sky130_fd_sc_hd__o211a_1 _1599_ (.A1(net23),
    .A2(_0772_),
    .B1(_0785_),
    .C1(_0727_),
    .X(_0802_));
 sky130_fd_sc_hd__and4_1 _1600_ (.A(net60),
    .B(net55),
    .C(net45),
    .D(net75),
    .X(_0803_));
 sky130_fd_sc_hd__or4_2 _1601_ (.A(net63),
    .B(net59),
    .C(net50),
    .D(net76),
    .X(_0804_));
 sky130_fd_sc_hd__nand2_1 _1602_ (.A(_0727_),
    .B(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__a31o_1 _1603_ (.A1(_0727_),
    .A2(_0785_),
    .A3(_0804_),
    .B1(net70),
    .X(_0806_));
 sky130_fd_sc_hd__o21ai_1 _1604_ (.A1(net73),
    .A2(_0802_),
    .B1(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__o211a_1 _1605_ (.A1(net73),
    .A2(_0802_),
    .B1(_0806_),
    .C1(_0787_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_1 _1606_ (.A(net33),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__nor2_1 _1607_ (.A(net94),
    .B(_0802_),
    .Y(_0810_));
 sky130_fd_sc_hd__nor2_1 _1608_ (.A(net69),
    .B(_0802_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _1609_ (.A(net44),
    .B(_0699_),
    .Y(_0812_));
 sky130_fd_sc_hd__or2_1 _1610_ (.A(net23),
    .B(net20),
    .X(_0813_));
 sky130_fd_sc_hd__a21oi_1 _1611_ (.A1(net26),
    .A2(_0812_),
    .B1(_0784_),
    .Y(_0814_));
 sky130_fd_sc_hd__nor2_1 _1612_ (.A(_0798_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__a211o_1 _1613_ (.A1(net26),
    .A2(_0771_),
    .B1(net17),
    .C1(_0700_),
    .X(_0816_));
 sky130_fd_sc_hd__o31a_1 _1614_ (.A1(_0811_),
    .A2(_0815_),
    .A3(_0816_),
    .B1(_0740_),
    .X(_0817_));
 sky130_fd_sc_hd__nor2_1 _1615_ (.A(_0691_),
    .B(_0726_),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _1616_ (.A(_0692_),
    .B(_0727_),
    .Y(_0819_));
 sky130_fd_sc_hd__or3_2 _1617_ (.A(_0691_),
    .B(net17),
    .C(_0803_),
    .X(_0820_));
 sky130_fd_sc_hd__a21o_1 _1618_ (.A1(net44),
    .A2(net76),
    .B1(net43),
    .X(_0821_));
 sky130_fd_sc_hd__and2_1 _1619_ (.A(net23),
    .B(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__a21o_2 _1620_ (.A1(net23),
    .A2(_0821_),
    .B1(net17),
    .X(_0823_));
 sky130_fd_sc_hd__or3_1 _1621_ (.A(_0723_),
    .B(_0798_),
    .C(_0823_),
    .X(_0824_));
 sky130_fd_sc_hd__o221a_1 _1622_ (.A1(net69),
    .A2(_0820_),
    .B1(_0823_),
    .B2(net112),
    .C1(net36),
    .X(_0825_));
 sky130_fd_sc_hd__a21o_1 _1623_ (.A1(net70),
    .A2(_0816_),
    .B1(_0820_),
    .X(_0826_));
 sky130_fd_sc_hd__a221o_1 _1624_ (.A1(_0824_),
    .A2(_0825_),
    .B1(_0826_),
    .B2(_0630_),
    .C1(net39),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_2 _1625_ (.A0(_0689_),
    .A1(_0709_),
    .S(net48),
    .X(_0828_));
 sky130_fd_sc_hd__mux2_2 _1626_ (.A0(net43),
    .A1(_0708_),
    .S(net48),
    .X(_0829_));
 sky130_fd_sc_hd__nand2_1 _1627_ (.A(net25),
    .B(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__a21o_1 _1628_ (.A1(net23),
    .A2(_0829_),
    .B1(_0726_),
    .X(_0831_));
 sky130_fd_sc_hd__nor2_2 _1629_ (.A(net98),
    .B(net105),
    .Y(_0832_));
 sky130_fd_sc_hd__nand2_2 _1630_ (.A(net100),
    .B(net112),
    .Y(_0833_));
 sky130_fd_sc_hd__nand2_2 _1631_ (.A(net102),
    .B(net93),
    .Y(_0834_));
 sky130_fd_sc_hd__nor2_2 _1632_ (.A(net98),
    .B(net69),
    .Y(_0835_));
 sky130_fd_sc_hd__nand2_1 _1633_ (.A(net101),
    .B(net71),
    .Y(_0836_));
 sky130_fd_sc_hd__o2111a_1 _1634_ (.A1(net20),
    .A2(net70),
    .B1(_0823_),
    .C1(net100),
    .D1(net85),
    .X(_0837_));
 sky130_fd_sc_hd__a211o_1 _1635_ (.A1(net48),
    .A2(_0708_),
    .B1(net64),
    .C1(net58),
    .X(_0838_));
 sky130_fd_sc_hd__nand2_1 _1636_ (.A(net53),
    .B(_0752_),
    .Y(_0839_));
 sky130_fd_sc_hd__a31o_2 _1637_ (.A1(net26),
    .A2(_0789_),
    .A3(_0839_),
    .B1(net21),
    .X(_0840_));
 sky130_fd_sc_hd__a311oi_2 _1638_ (.A1(net27),
    .A2(_0789_),
    .A3(_0839_),
    .B1(net21),
    .C1(net34),
    .Y(_0841_));
 sky130_fd_sc_hd__nand2_1 _1639_ (.A(net106),
    .B(_0677_),
    .Y(_0842_));
 sky130_fd_sc_hd__a311o_1 _1640_ (.A1(_0740_),
    .A2(_0831_),
    .A3(_0842_),
    .B1(_0841_),
    .C1(net40),
    .X(_0843_));
 sky130_fd_sc_hd__nand2_2 _1641_ (.A(net82),
    .B(_0832_),
    .Y(_0844_));
 sky130_fd_sc_hd__inv_2 _1642_ (.A(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__a2111o_1 _1643_ (.A1(net61),
    .A2(net56),
    .B1(net53),
    .C1(net79),
    .D1(net91),
    .X(_0846_));
 sky130_fd_sc_hd__o31a_2 _1644_ (.A1(net27),
    .A2(net94),
    .A3(_0828_),
    .B1(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__nand2_1 _1645_ (.A(net17),
    .B(_0772_),
    .Y(_0848_));
 sky130_fd_sc_hd__a21oi_1 _1646_ (.A1(_0847_),
    .A2(_0848_),
    .B1(_0844_),
    .Y(_0849_));
 sky130_fd_sc_hd__nor2_4 _1647_ (.A(net98),
    .B(net112),
    .Y(_0850_));
 sky130_fd_sc_hd__nand2_4 _1648_ (.A(net100),
    .B(net105),
    .Y(_0851_));
 sky130_fd_sc_hd__nor2_1 _1649_ (.A(net87),
    .B(_0851_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand2_2 _1650_ (.A(net83),
    .B(_0850_),
    .Y(_0853_));
 sky130_fd_sc_hd__and3_1 _1651_ (.A(_0654_),
    .B(_0656_),
    .C(net90),
    .X(_0854_));
 sky130_fd_sc_hd__nand2_1 _1652_ (.A(net27),
    .B(net90),
    .Y(_0855_));
 sky130_fd_sc_hd__a311o_1 _1653_ (.A1(net26),
    .A2(_0789_),
    .A3(_0839_),
    .B1(_0854_),
    .C1(_0667_),
    .X(_0856_));
 sky130_fd_sc_hd__a21oi_1 _1654_ (.A1(_0848_),
    .A2(_0856_),
    .B1(_0853_),
    .Y(_0857_));
 sky130_fd_sc_hd__o41a_1 _1655_ (.A1(_0837_),
    .A2(_0843_),
    .A3(_0849_),
    .A4(_0857_),
    .B1(net16),
    .X(_0858_));
 sky130_fd_sc_hd__o31a_1 _1656_ (.A1(_0809_),
    .A2(_0817_),
    .A3(_0827_),
    .B1(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__o21a_1 _1657_ (.A1(_0801_),
    .A2(_0859_),
    .B1(net8),
    .X(_0860_));
 sky130_fd_sc_hd__nand2b_1 _1658_ (.A_N(\logo_left[0] ),
    .B(\pix_x[0] ),
    .Y(_0861_));
 sky130_fd_sc_hd__and2_1 _1659_ (.A(_0599_),
    .B(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__nand2_2 _1660_ (.A(_0599_),
    .B(_0861_),
    .Y(_0863_));
 sky130_fd_sc_hd__a21oi_2 _1661_ (.A1(net62),
    .A2(net57),
    .B1(net93),
    .Y(_0864_));
 sky130_fd_sc_hd__nand2_2 _1662_ (.A(net24),
    .B(net96),
    .Y(_0865_));
 sky130_fd_sc_hd__nor2_1 _1663_ (.A(_0668_),
    .B(_0761_),
    .Y(_0866_));
 sky130_fd_sc_hd__a21oi_4 _1664_ (.A1(net21),
    .A2(_0762_),
    .B1(_0747_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand2_1 _1665_ (.A(net27),
    .B(net20),
    .Y(_0868_));
 sky130_fd_sc_hd__a21o_1 _1666_ (.A1(net19),
    .A2(_0742_),
    .B1(net102),
    .X(_0869_));
 sky130_fd_sc_hd__o21a_1 _1667_ (.A1(net19),
    .A2(net93),
    .B1(_0742_),
    .X(_0870_));
 sky130_fd_sc_hd__o2111a_1 _1668_ (.A1(net110),
    .A2(_0870_),
    .B1(_0869_),
    .C1(_0867_),
    .D1(_0865_),
    .X(_0871_));
 sky130_fd_sc_hd__nor2_1 _1669_ (.A(net100),
    .B(net70),
    .Y(_0872_));
 sky130_fd_sc_hd__or2_2 _1670_ (.A(net100),
    .B(net70),
    .X(_0873_));
 sky130_fd_sc_hd__and2_2 _1671_ (.A(net19),
    .B(_0732_),
    .X(_0874_));
 sky130_fd_sc_hd__a21o_1 _1672_ (.A1(net20),
    .A2(_0732_),
    .B1(_0872_),
    .X(_0875_));
 sky130_fd_sc_hd__a211o_1 _1673_ (.A1(_0711_),
    .A2(_0732_),
    .B1(_0798_),
    .C1(net102),
    .X(_0876_));
 sky130_fd_sc_hd__a21o_1 _1674_ (.A1(_0875_),
    .A2(_0876_),
    .B1(net87),
    .X(_0877_));
 sky130_fd_sc_hd__nor2_2 _1675_ (.A(net87),
    .B(_0778_),
    .Y(_0878_));
 sky130_fd_sc_hd__nand2_4 _1676_ (.A(net84),
    .B(_0777_),
    .Y(_0879_));
 sky130_fd_sc_hd__a21o_1 _1677_ (.A1(_0711_),
    .A2(_0732_),
    .B1(net96),
    .X(_0880_));
 sky130_fd_sc_hd__a21o_1 _1678_ (.A1(_0767_),
    .A2(_0880_),
    .B1(_0879_),
    .X(_0881_));
 sky130_fd_sc_hd__o2111a_1 _1679_ (.A1(net84),
    .A2(_0871_),
    .B1(_0877_),
    .C1(_0881_),
    .D1(net41),
    .X(_0882_));
 sky130_fd_sc_hd__o211a_4 _1680_ (.A1(net46),
    .A2(net79),
    .B1(net61),
    .C1(net56),
    .X(_0883_));
 sky130_fd_sc_hd__a211o_2 _1681_ (.A1(net54),
    .A2(net77),
    .B1(net65),
    .C1(_0655_),
    .X(_0884_));
 sky130_fd_sc_hd__o21ai_1 _1682_ (.A1(_0770_),
    .A2(_0883_),
    .B1(net69),
    .Y(_0885_));
 sky130_fd_sc_hd__a21o_1 _1683_ (.A1(_0733_),
    .A2(_0734_),
    .B1(net92),
    .X(_0886_));
 sky130_fd_sc_hd__a22o_1 _1684_ (.A1(net62),
    .A2(net57),
    .B1(net48),
    .B2(_0709_),
    .X(_0887_));
 sky130_fd_sc_hd__o2111a_1 _1685_ (.A1(net109),
    .A2(_0886_),
    .B1(_0887_),
    .C1(_0884_),
    .D1(_0885_),
    .X(_0888_));
 sky130_fd_sc_hd__and2_2 _1686_ (.A(net22),
    .B(_0693_),
    .X(_0889_));
 sky130_fd_sc_hd__o22a_1 _1687_ (.A1(net93),
    .A2(_0748_),
    .B1(_0828_),
    .B2(net110),
    .X(_0890_));
 sky130_fd_sc_hd__a21o_1 _1688_ (.A1(_0889_),
    .A2(_0890_),
    .B1(net66),
    .X(_0891_));
 sky130_fd_sc_hd__a21o_2 _1689_ (.A1(net22),
    .A2(_0693_),
    .B1(_0829_),
    .X(_0892_));
 sky130_fd_sc_hd__o21a_1 _1690_ (.A1(net32),
    .A2(_0892_),
    .B1(net37),
    .X(_0893_));
 sky130_fd_sc_hd__o21a_1 _1691_ (.A1(net109),
    .A2(_0889_),
    .B1(_0695_),
    .X(_0894_));
 sky130_fd_sc_hd__o221a_1 _1692_ (.A1(net34),
    .A2(_0888_),
    .B1(_0894_),
    .B2(net31),
    .C1(_0891_),
    .X(_0895_));
 sky130_fd_sc_hd__a211o_1 _1693_ (.A1(_0893_),
    .A2(_0895_),
    .B1(net12),
    .C1(_0882_),
    .X(_0896_));
 sky130_fd_sc_hd__o211a_2 _1694_ (.A1(net63),
    .A2(net59),
    .B1(net47),
    .C1(_0752_),
    .X(_0897_));
 sky130_fd_sc_hd__a211o_2 _1695_ (.A1(net61),
    .A2(net56),
    .B1(net53),
    .C1(_0751_),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_1 _1696_ (.A(_0710_),
    .B(_0884_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_1 _1697_ (.A(_0711_),
    .B(_0883_),
    .Y(_0900_));
 sky130_fd_sc_hd__a21oi_4 _1698_ (.A1(_0711_),
    .A2(_0883_),
    .B1(_0897_),
    .Y(_0901_));
 sky130_fd_sc_hd__nor2_1 _1699_ (.A(net106),
    .B(_0901_),
    .Y(_0902_));
 sky130_fd_sc_hd__nand2_1 _1700_ (.A(_0763_),
    .B(_0883_),
    .Y(_0903_));
 sky130_fd_sc_hd__a21oi_2 _1701_ (.A1(_0763_),
    .A2(_0883_),
    .B1(_0897_),
    .Y(_0904_));
 sky130_fd_sc_hd__mux2_1 _1702_ (.A0(_0901_),
    .A1(_0904_),
    .S(net107),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_1 _1703_ (.A(net43),
    .B(_0838_),
    .Y(_0906_));
 sky130_fd_sc_hd__o211a_1 _1704_ (.A1(net64),
    .A2(net58),
    .B1(net90),
    .C1(_0751_),
    .X(_0907_));
 sky130_fd_sc_hd__or2_1 _1705_ (.A(_0770_),
    .B(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__a211o_1 _1706_ (.A1(net27),
    .A2(_0794_),
    .B1(_0907_),
    .C1(_0770_),
    .X(_0909_));
 sky130_fd_sc_hd__nand2_1 _1707_ (.A(net81),
    .B(net68),
    .Y(_0910_));
 sky130_fd_sc_hd__o221a_1 _1708_ (.A1(net31),
    .A2(_0904_),
    .B1(_0910_),
    .B2(_0867_),
    .C1(net37),
    .X(_0911_));
 sky130_fd_sc_hd__o32a_1 _1709_ (.A1(_0698_),
    .A2(_0752_),
    .A3(_0884_),
    .B1(_0909_),
    .B2(net108),
    .X(_0912_));
 sky130_fd_sc_hd__o22a_1 _1710_ (.A1(net33),
    .A2(_0905_),
    .B1(_0912_),
    .B2(net66),
    .X(_0913_));
 sky130_fd_sc_hd__nor2_1 _1711_ (.A(_0761_),
    .B(_0838_),
    .Y(_0914_));
 sky130_fd_sc_hd__nand2_1 _1712_ (.A(net26),
    .B(_0790_),
    .Y(_0915_));
 sky130_fd_sc_hd__a211o_1 _1713_ (.A1(net27),
    .A2(_0790_),
    .B1(net21),
    .C1(net81),
    .X(_0916_));
 sky130_fd_sc_hd__o21a_1 _1714_ (.A1(net85),
    .A2(_0901_),
    .B1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__nand2_1 _1715_ (.A(net69),
    .B(_0897_),
    .Y(_0918_));
 sky130_fd_sc_hd__nor2_1 _1716_ (.A(net50),
    .B(net30),
    .Y(_0919_));
 sky130_fd_sc_hd__a211o_2 _1717_ (.A1(net60),
    .A2(net55),
    .B1(net50),
    .C1(net30),
    .X(_0920_));
 sky130_fd_sc_hd__a31o_1 _1718_ (.A1(_0900_),
    .A2(_0918_),
    .A3(_0920_),
    .B1(net66),
    .X(_0921_));
 sky130_fd_sc_hd__o221a_1 _1719_ (.A1(net33),
    .A2(_0840_),
    .B1(_0916_),
    .B2(net70),
    .C1(net40),
    .X(_0922_));
 sky130_fd_sc_hd__o211a_1 _1720_ (.A1(net102),
    .A2(_0917_),
    .B1(_0921_),
    .C1(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__a211o_1 _1721_ (.A1(_0911_),
    .A2(_0913_),
    .B1(_0923_),
    .C1(net16),
    .X(_0924_));
 sky130_fd_sc_hd__a21oi_1 _1722_ (.A1(_0896_),
    .A2(_0924_),
    .B1(net8),
    .Y(_0925_));
 sky130_fd_sc_hd__or3_1 _1723_ (.A(_0860_),
    .B(_0862_),
    .C(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__or3_1 _1724_ (.A(_0724_),
    .B(_0728_),
    .C(_0798_),
    .X(_0927_));
 sky130_fd_sc_hd__or3_1 _1725_ (.A(net97),
    .B(_0724_),
    .C(_0728_),
    .X(_0928_));
 sky130_fd_sc_hd__a21oi_1 _1726_ (.A1(_0736_),
    .A2(_0927_),
    .B1(net99),
    .Y(_0929_));
 sky130_fd_sc_hd__a41o_1 _1727_ (.A1(_0736_),
    .A2(_0744_),
    .A3(_0927_),
    .A4(_0928_),
    .B1(net99),
    .X(_0930_));
 sky130_fd_sc_hd__o2bb2a_1 _1728_ (.A1_N(net92),
    .A2_N(_0707_),
    .B1(_0673_),
    .B2(_0679_),
    .X(_0931_));
 sky130_fd_sc_hd__a31o_1 _1729_ (.A1(_0746_),
    .A2(_0930_),
    .A3(_0931_),
    .B1(net83),
    .X(_0932_));
 sky130_fd_sc_hd__a31o_1 _1730_ (.A1(net22),
    .A2(_0668_),
    .A3(net92),
    .B1(_0851_),
    .X(_0933_));
 sky130_fd_sc_hd__a21o_1 _1731_ (.A1(net97),
    .A2(_0718_),
    .B1(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__a211o_1 _1732_ (.A1(_0679_),
    .A2(net92),
    .B1(_0844_),
    .C1(_0673_),
    .X(_0935_));
 sky130_fd_sc_hd__o211a_1 _1733_ (.A1(net87),
    .A2(_0934_),
    .B1(_0935_),
    .C1(_0721_),
    .X(_0936_));
 sky130_fd_sc_hd__o2bb2a_1 _1734_ (.A1_N(_0700_),
    .A2_N(_0750_),
    .B1(_0733_),
    .B2(_0710_),
    .X(_0937_));
 sky130_fd_sc_hd__a221o_1 _1735_ (.A1(_0711_),
    .A2(_0732_),
    .B1(net30),
    .B2(_0700_),
    .C1(net92),
    .X(_0938_));
 sky130_fd_sc_hd__a21o_1 _1736_ (.A1(_0680_),
    .A2(_0766_),
    .B1(net95),
    .X(_0939_));
 sky130_fd_sc_hd__or2_1 _1737_ (.A(net95),
    .B(net18),
    .X(_0940_));
 sky130_fd_sc_hd__a21o_1 _1738_ (.A1(_0773_),
    .A2(_0915_),
    .B1(_0698_),
    .X(_0941_));
 sky130_fd_sc_hd__a211o_4 _1739_ (.A1(net46),
    .A2(_0675_),
    .B1(net63),
    .C1(net59),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _1740_ (.A0(net75),
    .A1(_0708_),
    .S(net50),
    .X(_0943_));
 sky130_fd_sc_hd__nor2_2 _1741_ (.A(_0761_),
    .B(_0942_),
    .Y(_0944_));
 sky130_fd_sc_hd__and3_2 _1742_ (.A(net24),
    .B(_0753_),
    .C(_0762_),
    .X(_0945_));
 sky130_fd_sc_hd__o21ai_1 _1743_ (.A1(_0944_),
    .A2(_0945_),
    .B1(net74),
    .Y(_0946_));
 sky130_fd_sc_hd__o21ai_4 _1744_ (.A1(_0761_),
    .A2(_0942_),
    .B1(_0785_),
    .Y(_0947_));
 sky130_fd_sc_hd__a21o_1 _1745_ (.A1(net23),
    .A2(_0790_),
    .B1(_0803_),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_1 _1746_ (.A(net74),
    .B(net72),
    .Y(_0949_));
 sky130_fd_sc_hd__nor2_2 _1747_ (.A(net81),
    .B(net68),
    .Y(_0950_));
 sky130_fd_sc_hd__nand2_4 _1748_ (.A(net85),
    .B(_0832_),
    .Y(_0951_));
 sky130_fd_sc_hd__mux2_1 _1749_ (.A0(_0718_),
    .A1(_0779_),
    .S(net95),
    .X(_0952_));
 sky130_fd_sc_hd__a31o_1 _1750_ (.A1(_0938_),
    .A2(_0939_),
    .A3(_0940_),
    .B1(net106),
    .X(_0953_));
 sky130_fd_sc_hd__a31o_1 _1751_ (.A1(_0941_),
    .A2(_0946_),
    .A3(_0953_),
    .B1(net67),
    .X(_0954_));
 sky130_fd_sc_hd__mux4_1 _1752_ (.A0(_0677_),
    .A1(_0790_),
    .A2(_0943_),
    .A3(_0783_),
    .S0(net24),
    .S1(net97),
    .X(_0955_));
 sky130_fd_sc_hd__nand2_1 _1753_ (.A(_0878_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__o211ai_1 _1754_ (.A1(_0745_),
    .A2(_0797_),
    .B1(_0948_),
    .C1(net35),
    .Y(_0957_));
 sky130_fd_sc_hd__o211a_1 _1755_ (.A1(_0951_),
    .A2(_0952_),
    .B1(_0956_),
    .C1(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__a32oi_4 _1756_ (.A1(_0781_),
    .A2(_0954_),
    .A3(_0958_),
    .B1(_0932_),
    .B2(_0936_),
    .Y(_0959_));
 sky130_fd_sc_hd__mux2_1 _1757_ (.A0(net77),
    .A1(_0752_),
    .S(net53),
    .X(_0960_));
 sky130_fd_sc_hd__nand2_2 _1758_ (.A(_0693_),
    .B(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__o22ai_2 _1759_ (.A1(net73),
    .A2(_0840_),
    .B1(_0961_),
    .B2(_0698_),
    .Y(_0962_));
 sky130_fd_sc_hd__or3b_1 _1760_ (.A(net46),
    .B(net91),
    .C_N(_0699_),
    .X(_0963_));
 sky130_fd_sc_hd__a31o_1 _1761_ (.A1(_0666_),
    .A2(net30),
    .A3(_0963_),
    .B1(net21),
    .X(_0964_));
 sky130_fd_sc_hd__nor2_1 _1762_ (.A(net105),
    .B(_0964_),
    .Y(_0965_));
 sky130_fd_sc_hd__o21a_1 _1763_ (.A1(_0962_),
    .A2(_0965_),
    .B1(_0630_),
    .X(_0966_));
 sky130_fd_sc_hd__or3_1 _1764_ (.A(_0818_),
    .B(net68),
    .C(_0897_),
    .X(_0967_));
 sky130_fd_sc_hd__a32o_1 _1765_ (.A1(_0819_),
    .A2(_0835_),
    .A3(_0898_),
    .B1(_0831_),
    .B2(net100),
    .X(_0968_));
 sky130_fd_sc_hd__and2_1 _1766_ (.A(net85),
    .B(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__nand2_1 _1767_ (.A(net85),
    .B(_0968_),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_2 _1768_ (.A(net82),
    .B(_0778_),
    .Y(_0971_));
 sky130_fd_sc_hd__nand2_4 _1769_ (.A(net89),
    .B(_0777_),
    .Y(_0972_));
 sky130_fd_sc_hd__a21o_1 _1770_ (.A1(_0666_),
    .A2(net30),
    .B1(net23),
    .X(_0973_));
 sky130_fd_sc_hd__nand2_1 _1771_ (.A(_0847_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__nor2_1 _1772_ (.A(net105),
    .B(net31),
    .Y(_0975_));
 sky130_fd_sc_hd__nand2_2 _1773_ (.A(net109),
    .B(_0740_),
    .Y(_0976_));
 sky130_fd_sc_hd__a221o_1 _1774_ (.A1(_0971_),
    .A2(_0974_),
    .B1(_0975_),
    .B2(_0831_),
    .C1(_0841_),
    .X(_0977_));
 sky130_fd_sc_hd__o31a_1 _1775_ (.A1(_0966_),
    .A2(_0969_),
    .A3(_0977_),
    .B1(net39),
    .X(_0978_));
 sky130_fd_sc_hd__o211a_1 _1776_ (.A1(net78),
    .A2(_0771_),
    .B1(net90),
    .C1(net26),
    .X(_0979_));
 sky130_fd_sc_hd__o32a_1 _1777_ (.A1(_0820_),
    .A2(net68),
    .A3(_0979_),
    .B1(_0851_),
    .B2(_0819_),
    .X(_0980_));
 sky130_fd_sc_hd__a211o_1 _1778_ (.A1(net90),
    .A2(_0820_),
    .B1(_0980_),
    .C1(net85),
    .X(_0981_));
 sky130_fd_sc_hd__or3_1 _1779_ (.A(net33),
    .B(_0807_),
    .C(_0947_),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _1780_ (.A1(_0797_),
    .A2(_0823_),
    .B1(_0918_),
    .B2(_0819_),
    .X(_0983_));
 sky130_fd_sc_hd__a211o_1 _1781_ (.A1(net90),
    .A2(_0823_),
    .B1(_0983_),
    .C1(net34),
    .X(_0984_));
 sky130_fd_sc_hd__a22o_2 _1782_ (.A1(net61),
    .A2(net56),
    .B1(net53),
    .B2(_0752_),
    .X(_0985_));
 sky130_fd_sc_hd__nand2_1 _1783_ (.A(_0727_),
    .B(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__a21o_1 _1784_ (.A1(net26),
    .A2(_0771_),
    .B1(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__nand2_1 _1785_ (.A(net90),
    .B(_0784_),
    .Y(_0988_));
 sky130_fd_sc_hd__o41a_1 _1786_ (.A1(net31),
    .A2(_0810_),
    .A3(_0815_),
    .A4(_0987_),
    .B1(net40),
    .X(_0989_));
 sky130_fd_sc_hd__a41o_1 _1787_ (.A1(_0981_),
    .A2(_0982_),
    .A3(_0984_),
    .A4(_0989_),
    .B1(net14),
    .X(_0990_));
 sky130_fd_sc_hd__o221a_1 _1788_ (.A1(net16),
    .A2(_0959_),
    .B1(_0978_),
    .B2(_0990_),
    .C1(net8),
    .X(_0991_));
 sky130_fd_sc_hd__o211ai_1 _1789_ (.A1(net110),
    .A2(_0886_),
    .B1(_0889_),
    .C1(_0885_),
    .Y(_0992_));
 sky130_fd_sc_hd__o21ai_1 _1790_ (.A1(_0873_),
    .A2(_0889_),
    .B1(net34),
    .Y(_0993_));
 sky130_fd_sc_hd__o21ai_1 _1791_ (.A1(_0829_),
    .A2(_0992_),
    .B1(_0993_),
    .Y(_0994_));
 sky130_fd_sc_hd__and4_1 _1792_ (.A(net37),
    .B(_0891_),
    .C(_0892_),
    .D(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__or2_1 _1793_ (.A(net93),
    .B(_0892_),
    .X(_0996_));
 sky130_fd_sc_hd__a31o_1 _1794_ (.A1(net19),
    .A2(_0732_),
    .A3(_0778_),
    .B1(net88),
    .X(_0997_));
 sky130_fd_sc_hd__a31o_1 _1795_ (.A1(_0777_),
    .A2(_0880_),
    .A3(_0996_),
    .B1(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__a21o_1 _1796_ (.A1(_0865_),
    .A2(_0867_),
    .B1(net33),
    .X(_0999_));
 sky130_fd_sc_hd__nor2_2 _1797_ (.A(net81),
    .B(_0851_),
    .Y(_1000_));
 sky130_fd_sc_hd__nand2_1 _1798_ (.A(net88),
    .B(_0850_),
    .Y(_1001_));
 sky130_fd_sc_hd__o221a_1 _1799_ (.A1(_0870_),
    .A2(_0976_),
    .B1(_1001_),
    .B2(_0742_),
    .C1(net41),
    .X(_1002_));
 sky130_fd_sc_hd__o2111a_1 _1800_ (.A1(_0874_),
    .A2(_0972_),
    .B1(_0998_),
    .C1(_0999_),
    .D1(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__o21ai_1 _1801_ (.A1(_0995_),
    .A2(_1003_),
    .B1(net15),
    .Y(_1004_));
 sky130_fd_sc_hd__o22a_1 _1802_ (.A1(_0710_),
    .A2(_0884_),
    .B1(_0898_),
    .B2(net91),
    .X(_1005_));
 sky130_fd_sc_hd__a21o_1 _1803_ (.A1(_0920_),
    .A2(_1005_),
    .B1(_0972_),
    .X(_1006_));
 sky130_fd_sc_hd__o21a_1 _1804_ (.A1(net86),
    .A2(_0901_),
    .B1(net40),
    .X(_1007_));
 sky130_fd_sc_hd__nand2_1 _1805_ (.A(net86),
    .B(_0778_),
    .Y(_1008_));
 sky130_fd_sc_hd__o211a_1 _1806_ (.A1(_0840_),
    .A2(_1008_),
    .B1(_1007_),
    .C1(_1006_),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _1807_ (.A1(net21),
    .A2(_0762_),
    .B1(_0883_),
    .B2(_0751_),
    .X(_1010_));
 sky130_fd_sc_hd__inv_2 _1808_ (.A(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__o221a_1 _1809_ (.A1(net32),
    .A2(_0901_),
    .B1(_1011_),
    .B2(net88),
    .C1(net37),
    .X(_1012_));
 sky130_fd_sc_hd__o32a_1 _1810_ (.A1(net31),
    .A2(_0798_),
    .A3(_0904_),
    .B1(_0976_),
    .B2(_0901_),
    .X(_1013_));
 sky130_fd_sc_hd__o211a_1 _1811_ (.A1(_0909_),
    .A2(_0972_),
    .B1(_1012_),
    .C1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__o21ai_1 _1812_ (.A1(_1009_),
    .A2(_1014_),
    .B1(net12),
    .Y(_1015_));
 sky130_fd_sc_hd__a311o_1 _1813_ (.A1(_0625_),
    .A2(_1004_),
    .A3(_1015_),
    .B1(_0863_),
    .C1(_0991_),
    .X(_1016_));
 sky130_fd_sc_hd__a21oi_1 _1814_ (.A1(_0926_),
    .A2(_1016_),
    .B1(_0602_),
    .Y(_1017_));
 sky130_fd_sc_hd__xnor2_2 _1815_ (.A(_0645_),
    .B(_0646_),
    .Y(_1018_));
 sky130_fd_sc_hd__inv_2 _1816_ (.A(_1018_),
    .Y(_1019_));
 sky130_fd_sc_hd__nor2_1 _1817_ (.A(net98),
    .B(_0808_),
    .Y(_1020_));
 sky130_fd_sc_hd__a21o_1 _1818_ (.A1(net98),
    .A2(_0816_),
    .B1(net81),
    .X(_1021_));
 sky130_fd_sc_hd__or3_1 _1819_ (.A(_0700_),
    .B(net17),
    .C(_0803_),
    .X(_1022_));
 sky130_fd_sc_hd__nor2_1 _1820_ (.A(net98),
    .B(net74),
    .Y(_1023_));
 sky130_fd_sc_hd__a21o_1 _1821_ (.A1(_1022_),
    .A2(_1023_),
    .B1(net85),
    .X(_1024_));
 sky130_fd_sc_hd__a21o_1 _1822_ (.A1(net26),
    .A2(_0786_),
    .B1(_0872_),
    .X(_1025_));
 sky130_fd_sc_hd__o32a_1 _1823_ (.A1(_0723_),
    .A2(_0823_),
    .A3(_0873_),
    .B1(_1025_),
    .B2(_0691_),
    .X(_1026_));
 sky130_fd_sc_hd__o22a_1 _1824_ (.A1(_1020_),
    .A2(_1021_),
    .B1(_1024_),
    .B2(_1026_),
    .X(_1027_));
 sky130_fd_sc_hd__a21oi_1 _1825_ (.A1(_0847_),
    .A2(_0848_),
    .B1(_0851_),
    .Y(_1028_));
 sky130_fd_sc_hd__and3_1 _1826_ (.A(_0711_),
    .B(_0823_),
    .C(_0832_),
    .X(_1029_));
 sky130_fd_sc_hd__a211o_1 _1827_ (.A1(net17),
    .A2(_0772_),
    .B1(net85),
    .C1(_0671_),
    .X(_1030_));
 sky130_fd_sc_hd__a32o_1 _1828_ (.A1(_0668_),
    .A2(_0872_),
    .A3(_0915_),
    .B1(_1030_),
    .B2(net66),
    .X(_1031_));
 sky130_fd_sc_hd__or3_1 _1829_ (.A(_1028_),
    .B(_1029_),
    .C(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _1830_ (.A(_0678_),
    .B(_0691_),
    .Y(_1033_));
 sky130_fd_sc_hd__nor2_1 _1831_ (.A(_0834_),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__a21o_1 _1832_ (.A1(_0727_),
    .A2(_0804_),
    .B1(_0919_),
    .X(_1035_));
 sky130_fd_sc_hd__o2111ai_1 _1833_ (.A1(net94),
    .A2(_0727_),
    .B1(_0950_),
    .C1(_1033_),
    .D1(_1035_),
    .Y(_1036_));
 sky130_fd_sc_hd__nand2_2 _1834_ (.A(net89),
    .B(net68),
    .Y(_1037_));
 sky130_fd_sc_hd__a211o_1 _1835_ (.A1(_0678_),
    .A2(_0831_),
    .B1(_1034_),
    .C1(_1037_),
    .X(_1038_));
 sky130_fd_sc_hd__a31o_1 _1836_ (.A1(_1032_),
    .A2(_1036_),
    .A3(_1038_),
    .B1(net40),
    .X(_1039_));
 sky130_fd_sc_hd__o211ai_1 _1837_ (.A1(net38),
    .A2(_1027_),
    .B1(_1039_),
    .C1(net16),
    .Y(_1040_));
 sky130_fd_sc_hd__nor2_1 _1838_ (.A(_0731_),
    .B(_0734_),
    .Y(_1041_));
 sky130_fd_sc_hd__o31ai_1 _1839_ (.A1(_0747_),
    .A2(_0755_),
    .A3(_1041_),
    .B1(_0740_),
    .Y(_1042_));
 sky130_fd_sc_hd__a21oi_1 _1840_ (.A1(_0735_),
    .A2(_0950_),
    .B1(net38),
    .Y(_1043_));
 sky130_fd_sc_hd__o311a_1 _1841_ (.A1(_0724_),
    .A2(_0728_),
    .A3(net32),
    .B1(_1042_),
    .C1(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__nand2_1 _1842_ (.A(net71),
    .B(_0755_),
    .Y(_1045_));
 sky130_fd_sc_hd__a2bb2o_1 _1843_ (.A1_N(_0702_),
    .A2_N(net69),
    .B1(_0797_),
    .B2(_0717_),
    .X(_1046_));
 sky130_fd_sc_hd__o21ba_1 _1844_ (.A1(net111),
    .A2(_0952_),
    .B1_N(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__or3b_1 _1845_ (.A(_0669_),
    .B(_0798_),
    .C_N(_0795_),
    .X(_1048_));
 sky130_fd_sc_hd__a31o_1 _1846_ (.A1(_0702_),
    .A2(_1045_),
    .A3(_1048_),
    .B1(net67),
    .X(_1049_));
 sky130_fd_sc_hd__o211a_1 _1847_ (.A1(net34),
    .A2(_1047_),
    .B1(_1049_),
    .C1(_1044_),
    .X(_1050_));
 sky130_fd_sc_hd__a21o_1 _1848_ (.A1(net24),
    .A2(_0943_),
    .B1(_0662_),
    .X(_1051_));
 sky130_fd_sc_hd__o221a_1 _1849_ (.A1(_0662_),
    .A2(_0945_),
    .B1(_1051_),
    .B2(net95),
    .C1(_0852_),
    .X(_1052_));
 sky130_fd_sc_hd__a21bo_1 _1850_ (.A1(_0680_),
    .A2(_0766_),
    .B1_N(net30),
    .X(_1053_));
 sky130_fd_sc_hd__nand2_1 _1851_ (.A(net22),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__a31o_1 _1852_ (.A1(_0630_),
    .A2(_0797_),
    .A3(_1051_),
    .B1(net42),
    .X(_1055_));
 sky130_fd_sc_hd__a311o_1 _1853_ (.A1(_0630_),
    .A2(net71),
    .A3(_1054_),
    .B1(_1055_),
    .C1(_1052_),
    .X(_1056_));
 sky130_fd_sc_hd__or3b_1 _1854_ (.A(_0662_),
    .B(net92),
    .C_N(_0791_),
    .X(_1057_));
 sky130_fd_sc_hd__o31a_1 _1855_ (.A1(_0662_),
    .A2(net95),
    .A3(_0945_),
    .B1(net111),
    .X(_1058_));
 sky130_fd_sc_hd__and3_1 _1856_ (.A(net35),
    .B(_1057_),
    .C(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__nor2_1 _1857_ (.A(_1056_),
    .B(_1059_),
    .Y(_1060_));
 sky130_fd_sc_hd__o21ai_1 _1858_ (.A1(net95),
    .A2(_0779_),
    .B1(net18),
    .Y(_1061_));
 sky130_fd_sc_hd__o21ai_1 _1859_ (.A1(_0777_),
    .A2(_0779_),
    .B1(_1053_),
    .Y(_1062_));
 sky130_fd_sc_hd__o21a_1 _1860_ (.A1(_1061_),
    .A2(_1062_),
    .B1(net87),
    .X(_1063_));
 sky130_fd_sc_hd__a2111oi_1 _1861_ (.A1(net35),
    .A2(_0793_),
    .B1(_1056_),
    .C1(_1059_),
    .D1(_1063_),
    .Y(_1064_));
 sky130_fd_sc_hd__o31a_1 _1862_ (.A1(net15),
    .A2(_1050_),
    .A3(net7),
    .B1(net8),
    .X(_1065_));
 sky130_fd_sc_hd__nor2_1 _1863_ (.A(_0732_),
    .B(_0770_),
    .Y(_1066_));
 sky130_fd_sc_hd__a31o_1 _1864_ (.A1(net110),
    .A2(_0884_),
    .A3(_0887_),
    .B1(net34),
    .X(_1067_));
 sky130_fd_sc_hd__a31o_1 _1865_ (.A1(net107),
    .A2(_0886_),
    .A3(_1066_),
    .B1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__or2_1 _1866_ (.A(net73),
    .B(_0887_),
    .X(_1069_));
 sky130_fd_sc_hd__a31o_1 _1867_ (.A1(_0748_),
    .A2(_0889_),
    .A3(_1069_),
    .B1(net66),
    .X(_1070_));
 sky130_fd_sc_hd__o21a_1 _1868_ (.A1(net107),
    .A2(_0767_),
    .B1(net38),
    .X(_1071_));
 sky130_fd_sc_hd__o211a_1 _1869_ (.A1(net73),
    .A2(_0693_),
    .B1(_0694_),
    .C1(_0663_),
    .X(_1072_));
 sky130_fd_sc_hd__or2_1 _1870_ (.A(net101),
    .B(_1072_),
    .X(_1073_));
 sky130_fd_sc_hd__and4_1 _1871_ (.A(_1068_),
    .B(_1070_),
    .C(_1071_),
    .D(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__o221a_1 _1872_ (.A1(net73),
    .A2(_0695_),
    .B1(net71),
    .B2(_0892_),
    .C1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__nand2_4 _1873_ (.A(net111),
    .B(net35),
    .Y(_1076_));
 sky130_fd_sc_hd__a21o_1 _1874_ (.A1(_0711_),
    .A2(_0732_),
    .B1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__and3_1 _1875_ (.A(net41),
    .B(_0881_),
    .C(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__a21o_1 _1876_ (.A1(net20),
    .A2(_0742_),
    .B1(net110),
    .X(_1079_));
 sky130_fd_sc_hd__a41o_1 _1877_ (.A1(_0865_),
    .A2(_0867_),
    .A3(_0869_),
    .A4(_1079_),
    .B1(net84),
    .X(_1080_));
 sky130_fd_sc_hd__a21o_1 _1878_ (.A1(net20),
    .A2(_0742_),
    .B1(_0844_),
    .X(_1081_));
 sky130_fd_sc_hd__o2111a_1 _1879_ (.A1(_0853_),
    .A2(_0874_),
    .B1(_1078_),
    .C1(_1080_),
    .D1(_1081_),
    .X(_1082_));
 sky130_fd_sc_hd__and3_1 _1880_ (.A(_0852_),
    .B(_0920_),
    .C(_1005_),
    .X(_1083_));
 sky130_fd_sc_hd__o21a_1 _1881_ (.A1(net21),
    .A2(_0914_),
    .B1(_0910_),
    .X(_1084_));
 sky130_fd_sc_hd__or3_1 _1882_ (.A(_0742_),
    .B(_0853_),
    .C(_0908_),
    .X(_1085_));
 sky130_fd_sc_hd__nand2_1 _1883_ (.A(_0910_),
    .B(_1008_),
    .Y(_1086_));
 sky130_fd_sc_hd__a211o_1 _1884_ (.A1(_0898_),
    .A2(_0942_),
    .B1(_1086_),
    .C1(net17),
    .X(_1087_));
 sky130_fd_sc_hd__o221a_1 _1885_ (.A1(net34),
    .A2(_0867_),
    .B1(_0904_),
    .B2(_1008_),
    .C1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__and3_1 _1886_ (.A(net37),
    .B(_1085_),
    .C(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__a211o_1 _1887_ (.A1(net36),
    .A2(_0905_),
    .B1(_1083_),
    .C1(_1084_),
    .X(_1090_));
 sky130_fd_sc_hd__a211o_1 _1888_ (.A1(_0705_),
    .A2(_1090_),
    .B1(_1089_),
    .C1(net15),
    .X(_1091_));
 sky130_fd_sc_hd__o311a_1 _1889_ (.A1(net12),
    .A2(_1075_),
    .A3(_1082_),
    .B1(_1091_),
    .C1(_0625_),
    .X(_1092_));
 sky130_fd_sc_hd__a211o_1 _1890_ (.A1(_1040_),
    .A2(_1065_),
    .B1(_1092_),
    .C1(_0863_),
    .X(_1093_));
 sky130_fd_sc_hd__nand2_1 _1891_ (.A(net91),
    .B(_0699_),
    .Y(_1094_));
 sky130_fd_sc_hd__o21a_1 _1892_ (.A1(net95),
    .A2(_0812_),
    .B1(net106),
    .X(_1095_));
 sky130_fd_sc_hd__o211a_1 _1893_ (.A1(net28),
    .A2(_0714_),
    .B1(net22),
    .C1(net111),
    .X(_1096_));
 sky130_fd_sc_hd__a311o_1 _1894_ (.A1(net22),
    .A2(_1053_),
    .A3(_1095_),
    .B1(_1096_),
    .C1(net101),
    .X(_1097_));
 sky130_fd_sc_hd__o211a_1 _1895_ (.A1(net28),
    .A2(_0714_),
    .B1(net74),
    .C1(net22),
    .X(_1098_));
 sky130_fd_sc_hd__a211o_1 _1896_ (.A1(net73),
    .A2(_0779_),
    .B1(_1098_),
    .C1(net99),
    .X(_1099_));
 sky130_fd_sc_hd__a21o_1 _1897_ (.A1(_1097_),
    .A2(_1099_),
    .B1(net84),
    .X(_1100_));
 sky130_fd_sc_hd__o21ai_1 _1898_ (.A1(_0700_),
    .A2(_0790_),
    .B1(net95),
    .Y(_1101_));
 sky130_fd_sc_hd__a31o_1 _1899_ (.A1(net22),
    .A2(_0791_),
    .A3(_1101_),
    .B1(_0879_),
    .X(_1102_));
 sky130_fd_sc_hd__or2_2 _1900_ (.A(net28),
    .B(_0812_),
    .X(_1103_));
 sky130_fd_sc_hd__o211a_1 _1901_ (.A1(net92),
    .A2(_0779_),
    .B1(_1103_),
    .C1(_0767_),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _1902_ (.A1(net71),
    .A2(_0755_),
    .B1(_0795_),
    .B2(_0670_),
    .X(_1105_));
 sky130_fd_sc_hd__o2bb2a_1 _1903_ (.A1_N(_0630_),
    .A2_N(_1105_),
    .B1(_0879_),
    .B2(_1104_),
    .X(_1106_));
 sky130_fd_sc_hd__o211a_1 _1904_ (.A1(_0702_),
    .A2(_1076_),
    .B1(_1106_),
    .C1(_1044_),
    .X(_1107_));
 sky130_fd_sc_hd__a311o_1 _1905_ (.A1(_1060_),
    .A2(_1100_),
    .A3(_1102_),
    .B1(_1107_),
    .C1(net15),
    .X(_1108_));
 sky130_fd_sc_hd__o22a_1 _1906_ (.A1(_0697_),
    .A2(_0847_),
    .B1(_0868_),
    .B2(_0771_),
    .X(_1109_));
 sky130_fd_sc_hd__or2_1 _1907_ (.A(net34),
    .B(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__a2111o_1 _1908_ (.A1(_0672_),
    .A2(net90),
    .B1(_0879_),
    .C1(_0914_),
    .D1(_0667_),
    .X(_1111_));
 sky130_fd_sc_hd__o41a_1 _1909_ (.A1(net66),
    .A2(_0677_),
    .A3(_0699_),
    .A4(_0765_),
    .B1(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__mux2_1 _1910_ (.A0(_0830_),
    .A1(_1033_),
    .S(_1023_),
    .X(_1113_));
 sky130_fd_sc_hd__a21o_1 _1911_ (.A1(_1035_),
    .A2(_1113_),
    .B1(net82),
    .X(_1114_));
 sky130_fd_sc_hd__and4_1 _1912_ (.A(net38),
    .B(_1110_),
    .C(_1112_),
    .D(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__nor2_2 _1913_ (.A(net101),
    .B(net73),
    .Y(_1116_));
 sky130_fd_sc_hd__o21a_1 _1914_ (.A1(net17),
    .A2(_0803_),
    .B1(net30),
    .X(_1117_));
 sky130_fd_sc_hd__o32a_1 _1915_ (.A1(_0822_),
    .A2(_0873_),
    .A3(_1117_),
    .B1(_1025_),
    .B2(_0700_),
    .X(_1118_));
 sky130_fd_sc_hd__a211o_1 _1916_ (.A1(_0728_),
    .A2(_1116_),
    .B1(_1118_),
    .C1(_1024_),
    .X(_1119_));
 sky130_fd_sc_hd__a22o_1 _1917_ (.A1(_0788_),
    .A2(_0832_),
    .B1(_0850_),
    .B2(_1022_),
    .X(_1120_));
 sky130_fd_sc_hd__o21ai_1 _1918_ (.A1(_1021_),
    .A2(_1120_),
    .B1(_1119_),
    .Y(_1121_));
 sky130_fd_sc_hd__a211o_1 _1919_ (.A1(net40),
    .A2(_1121_),
    .B1(_1115_),
    .C1(net13),
    .X(_1122_));
 sky130_fd_sc_hd__or2_1 _1920_ (.A(net109),
    .B(_0695_),
    .X(_1123_));
 sky130_fd_sc_hd__nand2_1 _1921_ (.A(net74),
    .B(_0919_),
    .Y(_1124_));
 sky130_fd_sc_hd__a31o_1 _1922_ (.A1(net20),
    .A2(_0742_),
    .A3(_1124_),
    .B1(net66),
    .X(_1125_));
 sky130_fd_sc_hd__nand2_1 _1923_ (.A(net23),
    .B(_0834_),
    .Y(_1126_));
 sky130_fd_sc_hd__a41o_1 _1924_ (.A1(_0813_),
    .A2(_0867_),
    .A3(_1079_),
    .A4(_1126_),
    .B1(net83),
    .X(_1127_));
 sky130_fd_sc_hd__and2_1 _1925_ (.A(_1125_),
    .B(_1127_),
    .X(_1128_));
 sky130_fd_sc_hd__a22o_1 _1926_ (.A1(_1074_),
    .A2(_1123_),
    .B1(_1128_),
    .B2(_1078_),
    .X(_1129_));
 sky130_fd_sc_hd__or3_1 _1927_ (.A(_0742_),
    .B(_0908_),
    .C(_1076_),
    .X(_1130_));
 sky130_fd_sc_hd__a221o_1 _1928_ (.A1(_0898_),
    .A2(_0942_),
    .B1(_1037_),
    .B2(net66),
    .C1(net17),
    .X(_1131_));
 sky130_fd_sc_hd__o221a_1 _1929_ (.A1(_0867_),
    .A2(_0879_),
    .B1(_0904_),
    .B2(_0951_),
    .C1(_1130_),
    .X(_1132_));
 sky130_fd_sc_hd__a31o_1 _1930_ (.A1(_0903_),
    .A2(_0918_),
    .A3(_0920_),
    .B1(net34),
    .X(_1133_));
 sky130_fd_sc_hd__a21o_1 _1931_ (.A1(_0732_),
    .A2(_0763_),
    .B1(_0671_),
    .X(_1134_));
 sky130_fd_sc_hd__nand2_1 _1932_ (.A(_0630_),
    .B(_1134_),
    .Y(_1135_));
 sky130_fd_sc_hd__a41o_1 _1933_ (.A1(net40),
    .A2(_0916_),
    .A3(_1133_),
    .A4(_1135_),
    .B1(net16),
    .X(_1136_));
 sky130_fd_sc_hd__a31o_1 _1934_ (.A1(net37),
    .A2(_1131_),
    .A3(_1132_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__o211a_1 _1935_ (.A1(net12),
    .A2(_1129_),
    .B1(_1137_),
    .C1(_0625_),
    .X(_1138_));
 sky130_fd_sc_hd__a311o_1 _1936_ (.A1(net8),
    .A2(_1108_),
    .A3(_1122_),
    .B1(_1138_),
    .C1(_0862_),
    .X(_1139_));
 sky130_fd_sc_hd__a31o_1 _1937_ (.A1(_0602_),
    .A2(_1093_),
    .A3(_1139_),
    .B1(_1018_),
    .X(_1140_));
 sky130_fd_sc_hd__nand2_1 _1938_ (.A(net111),
    .B(_0717_),
    .Y(_1141_));
 sky130_fd_sc_hd__a21o_1 _1939_ (.A1(_0725_),
    .A2(_0892_),
    .B1(net96),
    .X(_1142_));
 sky130_fd_sc_hd__a31o_1 _1940_ (.A1(_0768_),
    .A2(_1141_),
    .A3(_1142_),
    .B1(net32),
    .X(_1143_));
 sky130_fd_sc_hd__nor2_1 _1941_ (.A(_0866_),
    .B(_1061_),
    .Y(_1144_));
 sky130_fd_sc_hd__a21oi_1 _1942_ (.A1(net28),
    .A2(_0790_),
    .B1(_0765_),
    .Y(_1145_));
 sky130_fd_sc_hd__a21o_1 _1943_ (.A1(_0898_),
    .A2(_1145_),
    .B1(net95),
    .X(_1146_));
 sky130_fd_sc_hd__a31o_1 _1944_ (.A1(_0767_),
    .A2(_1103_),
    .A3(_1146_),
    .B1(_0853_),
    .X(_1147_));
 sky130_fd_sc_hd__a211o_1 _1945_ (.A1(net28),
    .A2(_0790_),
    .B1(_0765_),
    .C1(_0724_),
    .X(_1148_));
 sky130_fd_sc_hd__nor2_1 _1946_ (.A(net92),
    .B(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__and2_1 _1947_ (.A(net92),
    .B(_0768_),
    .X(_1150_));
 sky130_fd_sc_hd__or3_1 _1948_ (.A(_0976_),
    .B(_1149_),
    .C(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__nand2_1 _1949_ (.A(_0790_),
    .B(_0854_),
    .Y(_1152_));
 sky130_fd_sc_hd__a211o_1 _1950_ (.A1(_0668_),
    .A2(_0838_),
    .B1(_0761_),
    .C1(net96),
    .X(_1153_));
 sky130_fd_sc_hd__a221o_1 _1951_ (.A1(_0845_),
    .A2(_0937_),
    .B1(_0971_),
    .B2(_1148_),
    .C1(net42),
    .X(_1154_));
 sky130_fd_sc_hd__a21bo_1 _1952_ (.A1(net96),
    .A2(_0947_),
    .B1_N(_1153_),
    .X(_1155_));
 sky130_fd_sc_hd__a21oi_1 _1953_ (.A1(_0878_),
    .A2(_1155_),
    .B1(_1154_),
    .Y(_1156_));
 sky130_fd_sc_hd__o211a_1 _1954_ (.A1(_1076_),
    .A2(_1144_),
    .B1(_1147_),
    .C1(_1151_),
    .X(_1157_));
 sky130_fd_sc_hd__and3_1 _1955_ (.A(_1143_),
    .B(_1156_),
    .C(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__o221a_1 _1956_ (.A1(net101),
    .A2(_0718_),
    .B1(net68),
    .B2(_0673_),
    .C1(net83),
    .X(_1159_));
 sky130_fd_sc_hd__nand2_1 _1957_ (.A(net101),
    .B(_0713_),
    .Y(_1160_));
 sky130_fd_sc_hd__a22o_1 _1958_ (.A1(_0680_),
    .A2(net71),
    .B1(_0797_),
    .B2(_0920_),
    .X(_1161_));
 sky130_fd_sc_hd__or3_1 _1959_ (.A(net111),
    .B(_0673_),
    .C(net92),
    .X(_1162_));
 sky130_fd_sc_hd__a32oi_1 _1960_ (.A1(_0670_),
    .A2(_0697_),
    .A3(_0920_),
    .B1(_1161_),
    .B2(_0743_),
    .Y(_1163_));
 sky130_fd_sc_hd__a31o_1 _1961_ (.A1(net87),
    .A2(_1162_),
    .A3(_1163_),
    .B1(_0737_),
    .X(_1164_));
 sky130_fd_sc_hd__a22o_1 _1962_ (.A1(_1159_),
    .A2(_1160_),
    .B1(_1164_),
    .B2(_0930_),
    .X(_1165_));
 sky130_fd_sc_hd__a21o_1 _1963_ (.A1(net42),
    .A2(_1165_),
    .B1(net15),
    .X(_1166_));
 sky130_fd_sc_hd__nand2_1 _1964_ (.A(_0850_),
    .B(_0974_),
    .Y(_1167_));
 sky130_fd_sc_hd__nand2_1 _1965_ (.A(net98),
    .B(_0965_),
    .Y(_1168_));
 sky130_fd_sc_hd__a31o_1 _1966_ (.A1(_0967_),
    .A2(_1167_),
    .A3(_1168_),
    .B1(net81),
    .X(_1169_));
 sky130_fd_sc_hd__nand2b_1 _1967_ (.A_N(_0961_),
    .B(_1008_),
    .Y(_1170_));
 sky130_fd_sc_hd__a21o_1 _1968_ (.A1(_0727_),
    .A2(_0754_),
    .B1(net90),
    .X(_1171_));
 sky130_fd_sc_hd__a21boi_1 _1969_ (.A1(net91),
    .A2(_0986_),
    .B1_N(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__o221a_1 _1970_ (.A1(_0818_),
    .A2(_0897_),
    .B1(_1172_),
    .B2(net105),
    .C1(net36),
    .X(_1173_));
 sky130_fd_sc_hd__o2111a_1 _1971_ (.A1(_0707_),
    .A2(_0942_),
    .B1(_0985_),
    .C1(_0988_),
    .D1(_1000_),
    .X(_1174_));
 sky130_fd_sc_hd__nand2_1 _1972_ (.A(_0942_),
    .B(_0985_),
    .Y(_1175_));
 sky130_fd_sc_hd__o221a_1 _1973_ (.A1(net73),
    .A2(_0748_),
    .B1(_0813_),
    .B2(_0698_),
    .C1(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__and3b_1 _1974_ (.A_N(_0728_),
    .B(_0785_),
    .C(_0804_),
    .X(_1177_));
 sky130_fd_sc_hd__a31o_1 _1975_ (.A1(net61),
    .A2(net56),
    .A3(net43),
    .B1(net106),
    .X(_1178_));
 sky130_fd_sc_hd__a21oi_1 _1976_ (.A1(_0942_),
    .A2(_0985_),
    .B1(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__a211oi_1 _1977_ (.A1(net105),
    .A2(_0986_),
    .B1(_1179_),
    .C1(net66),
    .Y(_1180_));
 sky130_fd_sc_hd__a2bb2o_1 _1978_ (.A1_N(net31),
    .A2_N(_1176_),
    .B1(_1177_),
    .B2(_0950_),
    .X(_1181_));
 sky130_fd_sc_hd__o41a_1 _1979_ (.A1(_1173_),
    .A2(_1174_),
    .A3(_1180_),
    .A4(_1181_),
    .B1(net40),
    .X(_1182_));
 sky130_fd_sc_hd__a311o_1 _1980_ (.A1(net39),
    .A2(_1169_),
    .A3(_1170_),
    .B1(_1182_),
    .C1(net14),
    .X(_1183_));
 sky130_fd_sc_hd__o211a_1 _1981_ (.A1(_1158_),
    .A2(_1166_),
    .B1(_1183_),
    .C1(net8),
    .X(_1184_));
 sky130_fd_sc_hd__o21ai_1 _1982_ (.A1(_0716_),
    .A2(_0992_),
    .B1(net35),
    .Y(_1185_));
 sky130_fd_sc_hd__o221a_1 _1983_ (.A1(net110),
    .A2(_0828_),
    .B1(_0887_),
    .B2(net93),
    .C1(_0889_),
    .X(_1186_));
 sky130_fd_sc_hd__a31o_1 _1984_ (.A1(net109),
    .A2(net49),
    .A3(_0708_),
    .B1(_0889_),
    .X(_1187_));
 sky130_fd_sc_hd__o22a_1 _1985_ (.A1(net67),
    .A2(_1186_),
    .B1(_1187_),
    .B2(_0741_),
    .X(_1188_));
 sky130_fd_sc_hd__o22a_1 _1986_ (.A1(_0798_),
    .A2(_0906_),
    .B1(_1011_),
    .B2(net69),
    .X(_1189_));
 sky130_fd_sc_hd__o22a_1 _1987_ (.A1(_0769_),
    .A2(_0836_),
    .B1(_0874_),
    .B2(_1116_),
    .X(_1190_));
 sky130_fd_sc_hd__and3_1 _1988_ (.A(net62),
    .B(net57),
    .C(_0709_),
    .X(_1191_));
 sky130_fd_sc_hd__and2_1 _1989_ (.A(_0722_),
    .B(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__or3_1 _1990_ (.A(net19),
    .B(_0687_),
    .C(_0741_),
    .X(_1193_));
 sky130_fd_sc_hd__a21o_1 _1991_ (.A1(_1192_),
    .A2(_1193_),
    .B1(_1037_),
    .X(_1194_));
 sky130_fd_sc_hd__o21a_1 _1992_ (.A1(net24),
    .A2(net19),
    .B1(_0694_),
    .X(_1195_));
 sky130_fd_sc_hd__o221a_1 _1993_ (.A1(net88),
    .A2(_1190_),
    .B1(_1195_),
    .B2(_0720_),
    .C1(_1194_),
    .X(_1196_));
 sky130_fd_sc_hd__o211a_1 _1994_ (.A1(net32),
    .A2(_1189_),
    .B1(_1196_),
    .C1(net41),
    .X(_1197_));
 sky130_fd_sc_hd__a311o_1 _1995_ (.A1(_0893_),
    .A2(_1185_),
    .A3(_1188_),
    .B1(_1197_),
    .C1(net12),
    .X(_1198_));
 sky130_fd_sc_hd__a22o_1 _1996_ (.A1(net21),
    .A2(_0762_),
    .B1(_0829_),
    .B2(net29),
    .X(_1199_));
 sky130_fd_sc_hd__o32a_1 _1997_ (.A1(_0668_),
    .A2(net93),
    .A3(_0761_),
    .B1(_0828_),
    .B2(net25),
    .X(_1200_));
 sky130_fd_sc_hd__or3_1 _1998_ (.A(net29),
    .B(_0676_),
    .C(_0714_),
    .X(_1201_));
 sky130_fd_sc_hd__nand2_1 _1999_ (.A(_1200_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__a21oi_1 _2000_ (.A1(_1200_),
    .A2(_1201_),
    .B1(net110),
    .Y(_1203_));
 sky130_fd_sc_hd__nor2_1 _2001_ (.A(_0902_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__a22o_1 _2002_ (.A1(_0833_),
    .A2(_1010_),
    .B1(_1199_),
    .B2(net109),
    .X(_1205_));
 sky130_fd_sc_hd__a221o_1 _2003_ (.A1(_0740_),
    .A2(_1199_),
    .B1(_1205_),
    .B2(net83),
    .C1(net41),
    .X(_1206_));
 sky130_fd_sc_hd__o21ba_1 _2004_ (.A1(net32),
    .A2(_1204_),
    .B1_N(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__mux2_1 _2005_ (.A0(_0672_),
    .A1(_0898_),
    .S(_0684_),
    .X(_1208_));
 sky130_fd_sc_hd__nand2_1 _2006_ (.A(_0714_),
    .B(_0742_),
    .Y(_1209_));
 sky130_fd_sc_hd__a21oi_1 _2007_ (.A1(_0693_),
    .A2(_0960_),
    .B1(net105),
    .Y(_1210_));
 sky130_fd_sc_hd__a31o_1 _2008_ (.A1(net105),
    .A2(_1208_),
    .A3(_1209_),
    .B1(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__a21o_1 _2009_ (.A1(net20),
    .A2(_0883_),
    .B1(_0897_),
    .X(_1212_));
 sky130_fd_sc_hd__o21ai_1 _2010_ (.A1(_0671_),
    .A2(net76),
    .B1(_1212_),
    .Y(_1213_));
 sky130_fd_sc_hd__or2_1 _2011_ (.A(net70),
    .B(_0901_),
    .X(_1214_));
 sky130_fd_sc_hd__a21o_1 _2012_ (.A1(_1213_),
    .A2(_1214_),
    .B1(net31),
    .X(_1215_));
 sky130_fd_sc_hd__o211a_1 _2013_ (.A1(net33),
    .A2(_1211_),
    .B1(_1215_),
    .C1(_1007_),
    .X(_1216_));
 sky130_fd_sc_hd__o311a_1 _2014_ (.A1(net15),
    .A2(_1207_),
    .A3(_1216_),
    .B1(_1198_),
    .C1(_0625_),
    .X(_1217_));
 sky130_fd_sc_hd__a31oi_1 _2015_ (.A1(_0938_),
    .A2(_0939_),
    .A3(_1152_),
    .B1(_0844_),
    .Y(_1218_));
 sky130_fd_sc_hd__nor2_1 _2016_ (.A(_0768_),
    .B(_0976_),
    .Y(_1219_));
 sky130_fd_sc_hd__a221o_1 _2017_ (.A1(net35),
    .A2(_0866_),
    .B1(_0878_),
    .B2(_0944_),
    .C1(net42),
    .X(_1220_));
 sky130_fd_sc_hd__nor2_1 _2018_ (.A(_0864_),
    .B(_1076_),
    .Y(_1221_));
 sky130_fd_sc_hd__a32o_1 _2019_ (.A1(net95),
    .A2(_0878_),
    .A3(_0947_),
    .B1(_0948_),
    .B2(_1221_),
    .X(_1222_));
 sky130_fd_sc_hd__or4_1 _2020_ (.A(_1218_),
    .B(_1219_),
    .C(_1220_),
    .D(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__o21ai_1 _2021_ (.A1(_0944_),
    .A2(_0945_),
    .B1(net96),
    .Y(_1224_));
 sky130_fd_sc_hd__a21o_1 _2022_ (.A1(_1146_),
    .A2(_1224_),
    .B1(_0853_),
    .X(_1225_));
 sky130_fd_sc_hd__o21a_1 _2023_ (.A1(net106),
    .A2(_0718_),
    .B1(_0779_),
    .X(_1226_));
 sky130_fd_sc_hd__o32a_1 _2024_ (.A1(_0972_),
    .A2(_1149_),
    .A3(_1150_),
    .B1(_1226_),
    .B2(net32),
    .X(_1227_));
 sky130_fd_sc_hd__and3b_1 _2025_ (.A_N(_1223_),
    .B(_1225_),
    .C(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__a22oi_1 _2026_ (.A1(_0670_),
    .A2(_0680_),
    .B1(_0698_),
    .B2(_1178_),
    .Y(_1229_));
 sky130_fd_sc_hd__a211o_1 _2027_ (.A1(_0673_),
    .A2(_0686_),
    .B1(_1229_),
    .C1(net101),
    .X(_1230_));
 sky130_fd_sc_hd__a32oi_1 _2028_ (.A1(net87),
    .A2(_0930_),
    .A3(_1230_),
    .B1(_1159_),
    .B2(_0934_),
    .Y(_1231_));
 sky130_fd_sc_hd__o21ai_1 _2029_ (.A1(net38),
    .A2(_1231_),
    .B1(net13),
    .Y(_1232_));
 sky130_fd_sc_hd__or3_1 _2030_ (.A(net74),
    .B(net70),
    .C(_1177_),
    .X(_1233_));
 sky130_fd_sc_hd__o21ai_1 _2031_ (.A1(_0707_),
    .A2(_0942_),
    .B1(_0785_),
    .Y(_1234_));
 sky130_fd_sc_hd__nand2_1 _2032_ (.A(net74),
    .B(_1234_),
    .Y(_1235_));
 sky130_fd_sc_hd__a21o_1 _2033_ (.A1(_1233_),
    .A2(_1235_),
    .B1(net33),
    .X(_1236_));
 sky130_fd_sc_hd__a221o_1 _2034_ (.A1(_0947_),
    .A2(_0950_),
    .B1(_0971_),
    .B2(_0987_),
    .C1(net39),
    .X(_1237_));
 sky130_fd_sc_hd__a22o_1 _2035_ (.A1(_0797_),
    .A2(_1175_),
    .B1(_1234_),
    .B2(net70),
    .X(_1238_));
 sky130_fd_sc_hd__o2111a_1 _2036_ (.A1(_0684_),
    .A2(_0985_),
    .B1(_0692_),
    .C1(net105),
    .D1(_0727_),
    .X(_1239_));
 sky130_fd_sc_hd__o211a_1 _2037_ (.A1(_0690_),
    .A2(_0855_),
    .B1(_0985_),
    .C1(_0727_),
    .X(_1240_));
 sky130_fd_sc_hd__a211o_1 _2038_ (.A1(net112),
    .A2(_1240_),
    .B1(_1239_),
    .C1(net66),
    .X(_1241_));
 sky130_fd_sc_hd__a22o_1 _2039_ (.A1(net36),
    .A2(_0983_),
    .B1(_1238_),
    .B2(_0740_),
    .X(_1242_));
 sky130_fd_sc_hd__and4bb_1 _2040_ (.A_N(_1237_),
    .B_N(_1242_),
    .C(_1241_),
    .D(_1236_),
    .X(_1243_));
 sky130_fd_sc_hd__nor2_1 _2041_ (.A(_0777_),
    .B(_0961_),
    .Y(_1244_));
 sky130_fd_sc_hd__o21ai_1 _2042_ (.A1(_0962_),
    .A2(_1244_),
    .B1(net81),
    .Y(_1245_));
 sky130_fd_sc_hd__o2bb2a_1 _2043_ (.A1_N(_0974_),
    .A2_N(_0975_),
    .B1(_0964_),
    .B2(_0972_),
    .X(_1246_));
 sky130_fd_sc_hd__a41o_1 _2044_ (.A1(net39),
    .A2(_0970_),
    .A3(_1245_),
    .A4(_1246_),
    .B1(net14),
    .X(_1247_));
 sky130_fd_sc_hd__o221a_1 _2045_ (.A1(_1228_),
    .A2(_1232_),
    .B1(_1243_),
    .B2(_1247_),
    .C1(net8),
    .X(_1248_));
 sky130_fd_sc_hd__o2111a_1 _2046_ (.A1(net67),
    .A2(_1186_),
    .B1(_0994_),
    .C1(_0892_),
    .D1(net39),
    .X(_1249_));
 sky130_fd_sc_hd__mux2_1 _2047_ (.A0(_0874_),
    .A1(_0892_),
    .S(_1116_),
    .X(_1250_));
 sky130_fd_sc_hd__o211a_1 _2048_ (.A1(net110),
    .A2(net19),
    .B1(_0722_),
    .C1(_0732_),
    .X(_1251_));
 sky130_fd_sc_hd__o22a_1 _2049_ (.A1(_0906_),
    .A2(_1001_),
    .B1(_1251_),
    .B2(net31),
    .X(_1252_));
 sky130_fd_sc_hd__o221a_1 _2050_ (.A1(_0738_),
    .A2(_1189_),
    .B1(_1250_),
    .B2(net88),
    .C1(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__a211o_1 _2051_ (.A1(net41),
    .A2(_1253_),
    .B1(_1249_),
    .C1(net12),
    .X(_1254_));
 sky130_fd_sc_hd__or3_1 _2052_ (.A(net112),
    .B(net91),
    .C(_0901_),
    .X(_1255_));
 sky130_fd_sc_hd__a221o_1 _2053_ (.A1(_0715_),
    .A2(net70),
    .B1(_1213_),
    .B2(_1255_),
    .C1(net31),
    .X(_1256_));
 sky130_fd_sc_hd__o211a_1 _2054_ (.A1(net33),
    .A2(_0840_),
    .B1(_1007_),
    .C1(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__nand2_1 _2055_ (.A(net106),
    .B(_1199_),
    .Y(_1258_));
 sky130_fd_sc_hd__a31o_1 _2056_ (.A1(_1103_),
    .A2(_1200_),
    .A3(_1258_),
    .B1(_0741_),
    .X(_1259_));
 sky130_fd_sc_hd__a211o_1 _2057_ (.A1(_1012_),
    .A2(_1259_),
    .B1(_1257_),
    .C1(net15),
    .X(_1260_));
 sky130_fd_sc_hd__a311o_1 _2058_ (.A1(_0625_),
    .A2(_1254_),
    .A3(_1260_),
    .B1(_0862_),
    .C1(_1248_),
    .X(_1261_));
 sky130_fd_sc_hd__o311a_1 _2059_ (.A1(_0863_),
    .A2(_1184_),
    .A3(_1217_),
    .B1(_1261_),
    .C1(_0602_),
    .X(_1262_));
 sky130_fd_sc_hd__a22o_1 _2060_ (.A1(_0762_),
    .A2(_0770_),
    .B1(_0960_),
    .B2(net29),
    .X(_1263_));
 sky130_fd_sc_hd__o31a_1 _2061_ (.A1(net25),
    .A2(_0828_),
    .A3(_0834_),
    .B1(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__o221a_1 _2062_ (.A1(net23),
    .A2(_0752_),
    .B1(_0786_),
    .B2(_0669_),
    .C1(_1094_),
    .X(_1265_));
 sky130_fd_sc_hd__o2bb2a_1 _2063_ (.A1_N(_0630_),
    .A2_N(_0961_),
    .B1(_1037_),
    .B2(_1264_),
    .X(_1266_));
 sky130_fd_sc_hd__o2bb2a_1 _2064_ (.A1_N(net36),
    .A2_N(_1211_),
    .B1(_1265_),
    .B2(_0951_),
    .X(_1267_));
 sky130_fd_sc_hd__a2111o_1 _2065_ (.A1(net46),
    .A2(_0675_),
    .B1(net79),
    .C1(net63),
    .D1(net59),
    .X(_1268_));
 sky130_fd_sc_hd__nand2_1 _2066_ (.A(_0985_),
    .B(_1268_),
    .Y(_1269_));
 sky130_fd_sc_hd__o31a_1 _2067_ (.A1(net86),
    .A2(_1179_),
    .A3(_1269_),
    .B1(net34),
    .X(_1270_));
 sky130_fd_sc_hd__a21oi_1 _2068_ (.A1(_0754_),
    .A2(_1268_),
    .B1(_0798_),
    .Y(_1271_));
 sky130_fd_sc_hd__a21o_1 _2069_ (.A1(net72),
    .A2(_1269_),
    .B1(_1271_),
    .X(_1272_));
 sky130_fd_sc_hd__a21oi_1 _2070_ (.A1(_0786_),
    .A2(_0864_),
    .B1(_0907_),
    .Y(_1273_));
 sky130_fd_sc_hd__a221o_1 _2071_ (.A1(net17),
    .A2(_0769_),
    .B1(_0786_),
    .B2(_0864_),
    .C1(_0907_),
    .X(_1274_));
 sky130_fd_sc_hd__a221o_1 _2072_ (.A1(net72),
    .A2(_1269_),
    .B1(_1274_),
    .B2(net108),
    .C1(_1271_),
    .X(_1275_));
 sky130_fd_sc_hd__nor2_1 _2073_ (.A(_0710_),
    .B(_0728_),
    .Y(_1276_));
 sky130_fd_sc_hd__a31oi_1 _2074_ (.A1(_0754_),
    .A2(_0950_),
    .A3(_1276_),
    .B1(net39),
    .Y(_1277_));
 sky130_fd_sc_hd__a22o_1 _2075_ (.A1(net27),
    .A2(_0794_),
    .B1(_0851_),
    .B2(_0687_),
    .X(_1278_));
 sky130_fd_sc_hd__a211o_1 _2076_ (.A1(net27),
    .A2(_0753_),
    .B1(net74),
    .C1(net100),
    .X(_1279_));
 sky130_fd_sc_hd__a221o_1 _2077_ (.A1(net25),
    .A2(_0839_),
    .B1(_1278_),
    .B2(_1279_),
    .C1(net82),
    .X(_1280_));
 sky130_fd_sc_hd__o211a_1 _2078_ (.A1(_1270_),
    .A2(_1275_),
    .B1(_1277_),
    .C1(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__a31o_1 _2079_ (.A1(net37),
    .A2(_1266_),
    .A3(_1267_),
    .B1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__o211ai_2 _2080_ (.A1(_0761_),
    .A2(_0838_),
    .B1(_0694_),
    .C1(_0725_),
    .Y(_1283_));
 sky130_fd_sc_hd__a22oi_1 _2081_ (.A1(_0949_),
    .A2(_1148_),
    .B1(_1283_),
    .B2(net72),
    .Y(_1284_));
 sky130_fd_sc_hd__nand2_1 _2082_ (.A(_1000_),
    .B(_1283_),
    .Y(_1285_));
 sky130_fd_sc_hd__o221a_1 _2083_ (.A1(net29),
    .A2(_0714_),
    .B1(_0865_),
    .B2(_0699_),
    .C1(_0915_),
    .X(_1286_));
 sky130_fd_sc_hd__or3_1 _2084_ (.A(net67),
    .B(_0798_),
    .C(_1103_),
    .X(_1287_));
 sky130_fd_sc_hd__nand2_1 _2085_ (.A(net96),
    .B(_1283_),
    .Y(_1288_));
 sky130_fd_sc_hd__a21o_1 _2086_ (.A1(_1142_),
    .A2(_1288_),
    .B1(_0951_),
    .X(_1289_));
 sky130_fd_sc_hd__a31o_1 _2087_ (.A1(_0767_),
    .A2(_1103_),
    .A3(_1152_),
    .B1(_0851_),
    .X(_1290_));
 sky130_fd_sc_hd__o221a_1 _2088_ (.A1(_0779_),
    .A2(_1076_),
    .B1(_1086_),
    .B2(_1145_),
    .C1(net38),
    .X(_1291_));
 sky130_fd_sc_hd__o211a_1 _2089_ (.A1(net89),
    .A2(_1290_),
    .B1(_1291_),
    .C1(_1287_),
    .X(_1292_));
 sky130_fd_sc_hd__o221a_1 _2090_ (.A1(net31),
    .A2(_1284_),
    .B1(_1286_),
    .B2(_0879_),
    .C1(_1285_),
    .X(_1293_));
 sky130_fd_sc_hd__and3_1 _2091_ (.A(_1289_),
    .B(_1292_),
    .C(_1293_),
    .X(_1294_));
 sky130_fd_sc_hd__a221o_1 _2092_ (.A1(net71),
    .A2(_0747_),
    .B1(_0920_),
    .B2(_0670_),
    .C1(net83),
    .X(_1295_));
 sky130_fd_sc_hd__o2bb2a_1 _2093_ (.A1_N(net32),
    .A2_N(_1295_),
    .B1(net68),
    .B2(_0728_),
    .X(_1296_));
 sky130_fd_sc_hd__o21a_1 _2094_ (.A1(_0673_),
    .A2(_0836_),
    .B1(net83),
    .X(_1297_));
 sky130_fd_sc_hd__a21o_1 _2095_ (.A1(_0725_),
    .A2(_0892_),
    .B1(net109),
    .X(_1298_));
 sky130_fd_sc_hd__nand2_1 _2096_ (.A(_0713_),
    .B(_0778_),
    .Y(_1299_));
 sky130_fd_sc_hd__a31o_1 _2097_ (.A1(_1297_),
    .A2(_1298_),
    .A3(_1299_),
    .B1(_1296_),
    .X(_1300_));
 sky130_fd_sc_hd__a22o_1 _2098_ (.A1(net75),
    .A2(_0835_),
    .B1(_0850_),
    .B2(_0743_),
    .X(_1301_));
 sky130_fd_sc_hd__nand2_1 _2099_ (.A(net87),
    .B(_1301_),
    .Y(_0101_));
 sky130_fd_sc_hd__a31o_1 _2100_ (.A1(net42),
    .A2(_1300_),
    .A3(_0101_),
    .B1(net15),
    .X(_0102_));
 sky130_fd_sc_hd__a2bb2o_1 _2101_ (.A1_N(_1294_),
    .A2_N(_0102_),
    .B1(net16),
    .B2(_1282_),
    .X(_0103_));
 sky130_fd_sc_hd__o21a_1 _2102_ (.A1(_0899_),
    .A2(_0945_),
    .B1(_0797_),
    .X(_0104_));
 sky130_fd_sc_hd__o21a_1 _2103_ (.A1(_1203_),
    .A2(_0104_),
    .B1(net35),
    .X(_0105_));
 sky130_fd_sc_hd__a21o_1 _2104_ (.A1(net19),
    .A2(_0883_),
    .B1(_0945_),
    .X(_0106_));
 sky130_fd_sc_hd__o211a_1 _2105_ (.A1(_0689_),
    .A2(_0836_),
    .B1(_1212_),
    .C1(net88),
    .X(_0107_));
 sky130_fd_sc_hd__a31o_1 _2106_ (.A1(net83),
    .A2(_0873_),
    .A3(_0106_),
    .B1(net37),
    .X(_0108_));
 sky130_fd_sc_hd__o311a_1 _2107_ (.A1(_0679_),
    .A2(_0765_),
    .A3(_0805_),
    .B1(_0878_),
    .C1(_0750_),
    .X(_0109_));
 sky130_fd_sc_hd__a211o_1 _2108_ (.A1(_0879_),
    .A2(_1199_),
    .B1(_0109_),
    .C1(net41),
    .X(_0110_));
 sky130_fd_sc_hd__o311a_1 _2109_ (.A1(_0105_),
    .A2(_0107_),
    .A3(_0108_),
    .B1(_0110_),
    .C1(net12),
    .X(_0111_));
 sky130_fd_sc_hd__and4bb_1 _2110_ (.A_N(_0662_),
    .B_N(_0716_),
    .C(_0693_),
    .D(net109),
    .X(_0112_));
 sky130_fd_sc_hd__a311o_1 _2111_ (.A1(net106),
    .A2(_0886_),
    .A3(_0928_),
    .B1(_0112_),
    .C1(_0720_),
    .X(_0113_));
 sky130_fd_sc_hd__o211a_1 _2112_ (.A1(_0663_),
    .A2(_0687_),
    .B1(_0693_),
    .C1(net18),
    .X(_0114_));
 sky130_fd_sc_hd__o211a_1 _2113_ (.A1(_0687_),
    .A2(_0748_),
    .B1(_0887_),
    .C1(_0663_),
    .X(_0115_));
 sky130_fd_sc_hd__o221a_1 _2114_ (.A1(net101),
    .A2(_0114_),
    .B1(_0115_),
    .B2(net67),
    .C1(net38),
    .X(_0116_));
 sky130_fd_sc_hd__nand2_1 _2115_ (.A(_0113_),
    .B(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__and2_1 _2116_ (.A(net109),
    .B(_1195_),
    .X(_0118_));
 sky130_fd_sc_hd__a31oi_1 _2117_ (.A1(net107),
    .A2(_0693_),
    .A3(net18),
    .B1(_0118_),
    .Y(_0119_));
 sky130_fd_sc_hd__a31o_1 _2118_ (.A1(net29),
    .A2(net19),
    .A3(_0709_),
    .B1(net107),
    .X(_0120_));
 sky130_fd_sc_hd__a21o_1 _2119_ (.A1(net19),
    .A2(_0883_),
    .B1(_0698_),
    .X(_0121_));
 sky130_fd_sc_hd__a21o_1 _2120_ (.A1(_0120_),
    .A2(_0121_),
    .B1(net102),
    .X(_0122_));
 sky130_fd_sc_hd__o31a_1 _2121_ (.A1(net109),
    .A2(net52),
    .A3(net77),
    .B1(net83),
    .X(_0123_));
 sky130_fd_sc_hd__a31o_1 _2122_ (.A1(_0722_),
    .A2(_1191_),
    .A3(_0123_),
    .B1(net35),
    .X(_0124_));
 sky130_fd_sc_hd__o21a_1 _2123_ (.A1(_0778_),
    .A2(_1195_),
    .B1(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__a22o_1 _2124_ (.A1(net25),
    .A2(_0835_),
    .B1(_1191_),
    .B2(_0722_),
    .X(_0126_));
 sky130_fd_sc_hd__and4_1 _2125_ (.A(net89),
    .B(_0725_),
    .C(_0766_),
    .D(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__a21oi_1 _2126_ (.A1(_0122_),
    .A2(_0125_),
    .B1(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__o221a_1 _2127_ (.A1(_0117_),
    .A2(_0119_),
    .B1(_0128_),
    .B2(net38),
    .C1(net15),
    .X(_0129_));
 sky130_fd_sc_hd__o21a_1 _2128_ (.A1(_0111_),
    .A2(_0129_),
    .B1(_0625_),
    .X(_0130_));
 sky130_fd_sc_hd__a211o_1 _2129_ (.A1(net8),
    .A2(_0103_),
    .B1(_0130_),
    .C1(_0863_),
    .X(_0131_));
 sky130_fd_sc_hd__a21oi_1 _2130_ (.A1(_1142_),
    .A2(_1288_),
    .B1(_0851_),
    .Y(_0132_));
 sky130_fd_sc_hd__a21oi_1 _2131_ (.A1(_0725_),
    .A2(_0892_),
    .B1(net68),
    .Y(_0133_));
 sky130_fd_sc_hd__a2111o_1 _2132_ (.A1(net99),
    .A2(_1148_),
    .B1(_0132_),
    .C1(_0133_),
    .D1(net84),
    .X(_0134_));
 sky130_fd_sc_hd__and3_1 _2133_ (.A(net106),
    .B(_1101_),
    .C(_1153_),
    .X(_0135_));
 sky130_fd_sc_hd__a211oi_1 _2134_ (.A1(net111),
    .A2(_0779_),
    .B1(_0135_),
    .C1(net101),
    .Y(_0136_));
 sky130_fd_sc_hd__nand2_1 _2135_ (.A(_0835_),
    .B(_0937_),
    .Y(_0137_));
 sky130_fd_sc_hd__o211ai_1 _2136_ (.A1(_0833_),
    .A2(_1145_),
    .B1(_0137_),
    .C1(net84),
    .Y(_0138_));
 sky130_fd_sc_hd__or3b_1 _2137_ (.A(_0138_),
    .B(_0136_),
    .C_N(_1290_),
    .X(_0139_));
 sky130_fd_sc_hd__o211a_1 _2138_ (.A1(net97),
    .A2(_0725_),
    .B1(_0743_),
    .C1(_0850_),
    .X(_0140_));
 sky130_fd_sc_hd__a211o_1 _2139_ (.A1(net32),
    .A2(_1295_),
    .B1(_0140_),
    .C1(_0929_),
    .X(_0141_));
 sky130_fd_sc_hd__a21oi_1 _2140_ (.A1(_0713_),
    .A2(_0873_),
    .B1(_0717_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _2141_ (.A(_1297_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__a31o_1 _2142_ (.A1(net42),
    .A2(_0141_),
    .A3(_0143_),
    .B1(net15),
    .X(_0144_));
 sky130_fd_sc_hd__a31o_1 _2143_ (.A1(net37),
    .A2(_0134_),
    .A3(_0139_),
    .B1(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__a21o_1 _2144_ (.A1(_0754_),
    .A2(_1268_),
    .B1(net94),
    .X(_0146_));
 sky130_fd_sc_hd__a21oi_1 _2145_ (.A1(_1171_),
    .A2(_0146_),
    .B1(_0778_),
    .Y(_0147_));
 sky130_fd_sc_hd__a211o_1 _2146_ (.A1(net98),
    .A2(_1272_),
    .B1(_0147_),
    .C1(_1270_),
    .X(_0148_));
 sky130_fd_sc_hd__and3_1 _2147_ (.A(net98),
    .B(_0813_),
    .C(_1176_),
    .X(_0149_));
 sky130_fd_sc_hd__o221a_1 _2148_ (.A1(_0829_),
    .A2(_0855_),
    .B1(_0942_),
    .B2(_0707_),
    .C1(_0985_),
    .X(_0150_));
 sky130_fd_sc_hd__nor2_1 _2149_ (.A(_0851_),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__a31o_1 _2150_ (.A1(_0754_),
    .A2(_0988_),
    .A3(_1276_),
    .B1(net68),
    .X(_0152_));
 sky130_fd_sc_hd__or4b_1 _2151_ (.A(net82),
    .B(_0149_),
    .C(_0151_),
    .D_N(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__and3_1 _2152_ (.A(_0950_),
    .B(_0973_),
    .C(_1273_),
    .X(_0154_));
 sky130_fd_sc_hd__a221o_1 _2153_ (.A1(net33),
    .A2(_0961_),
    .B1(_0964_),
    .B2(_1000_),
    .C1(net40),
    .X(_0155_));
 sky130_fd_sc_hd__nor2_1 _2154_ (.A(_0154_),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__a311o_1 _2155_ (.A1(net40),
    .A2(_0148_),
    .A3(_0153_),
    .B1(_0156_),
    .C1(net14),
    .X(_0157_));
 sky130_fd_sc_hd__o21a_1 _2156_ (.A1(_0899_),
    .A2(_0945_),
    .B1(net106),
    .X(_0158_));
 sky130_fd_sc_hd__o21a_1 _2157_ (.A1(_0902_),
    .A2(_0158_),
    .B1(net36),
    .X(_0159_));
 sky130_fd_sc_hd__a211o_1 _2158_ (.A1(_0711_),
    .A2(_0883_),
    .B1(_0897_),
    .C1(net72),
    .X(_0160_));
 sky130_fd_sc_hd__o211a_1 _2159_ (.A1(net69),
    .A2(_1212_),
    .B1(_0160_),
    .C1(_0630_),
    .X(_0161_));
 sky130_fd_sc_hd__a21oi_1 _2160_ (.A1(_1208_),
    .A2(_1209_),
    .B1(_0951_),
    .Y(_0162_));
 sky130_fd_sc_hd__o2111a_1 _2161_ (.A1(_0689_),
    .A2(_0834_),
    .B1(_1212_),
    .C1(net68),
    .D1(net86),
    .X(_0163_));
 sky130_fd_sc_hd__or4_1 _2162_ (.A(net37),
    .B(_0161_),
    .C(_0162_),
    .D(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__a31o_1 _2163_ (.A1(_0720_),
    .A2(_0951_),
    .A3(_1199_),
    .B1(net41),
    .X(_0165_));
 sky130_fd_sc_hd__a221o_1 _2164_ (.A1(net36),
    .A2(_1010_),
    .B1(_1202_),
    .B2(net88),
    .C1(_0165_),
    .X(_0166_));
 sky130_fd_sc_hd__o211a_1 _2165_ (.A1(net93),
    .A2(_0693_),
    .B1(_0892_),
    .C1(net107),
    .X(_0167_));
 sky130_fd_sc_hd__o211a_1 _2166_ (.A1(_0118_),
    .A2(_0167_),
    .B1(_0113_),
    .C1(_0116_),
    .X(_0168_));
 sky130_fd_sc_hd__o211a_1 _2167_ (.A1(net96),
    .A2(_0874_),
    .B1(_1195_),
    .C1(_0120_),
    .X(_0169_));
 sky130_fd_sc_hd__a211o_1 _2168_ (.A1(_0769_),
    .A2(_0874_),
    .B1(net67),
    .C1(net71),
    .X(_0170_));
 sky130_fd_sc_hd__o311a_1 _2169_ (.A1(net88),
    .A2(_0834_),
    .A3(_1192_),
    .B1(_0170_),
    .C1(net41),
    .X(_0171_));
 sky130_fd_sc_hd__and2b_1 _2170_ (.A_N(_0866_),
    .B(_0126_),
    .X(_0172_));
 sky130_fd_sc_hd__o22a_1 _2171_ (.A1(_0720_),
    .A2(_0169_),
    .B1(_0172_),
    .B2(net84),
    .X(_0173_));
 sky130_fd_sc_hd__o211ai_1 _2172_ (.A1(_0159_),
    .A2(_0164_),
    .B1(_0166_),
    .C1(net13),
    .Y(_0174_));
 sky130_fd_sc_hd__a221o_1 _2173_ (.A1(_0996_),
    .A2(_0168_),
    .B1(_0171_),
    .B2(_0173_),
    .C1(net12),
    .X(_0175_));
 sky130_fd_sc_hd__a21oi_1 _2174_ (.A1(_0174_),
    .A2(_0175_),
    .B1(net8),
    .Y(_0176_));
 sky130_fd_sc_hd__a311o_1 _2175_ (.A1(_0624_),
    .A2(_0145_),
    .A3(_0157_),
    .B1(_0176_),
    .C1(_0862_),
    .X(_0177_));
 sky130_fd_sc_hd__a21oi_1 _2176_ (.A1(_0131_),
    .A2(_0177_),
    .B1(_0602_),
    .Y(_0178_));
 sky130_fd_sc_hd__or3_2 _2177_ (.A(_1019_),
    .B(_1262_),
    .C(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__a21oi_1 _2178_ (.A1(_0605_),
    .A2(_0623_),
    .B1(_0603_),
    .Y(_0180_));
 sky130_fd_sc_hd__xor2_1 _2179_ (.A(\logo_top[9] ),
    .B(\pix_y[9] ),
    .X(_0181_));
 sky130_fd_sc_hd__a21o_1 _2180_ (.A1(_0519_),
    .A2(net118),
    .B1(_0181_),
    .X(_0182_));
 sky130_fd_sc_hd__and4_1 _2181_ (.A(net125),
    .B(_0533_),
    .C(_0180_),
    .D(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__nand2_1 _2182_ (.A(_0520_),
    .B(\pix_y[7] ),
    .Y(_0184_));
 sky130_fd_sc_hd__a21o_1 _2183_ (.A1(net125),
    .A2(_0533_),
    .B1(_0182_),
    .X(_0185_));
 sky130_fd_sc_hd__a21oi_1 _2184_ (.A1(_0180_),
    .A2(_0184_),
    .B1(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__or2_1 _2185_ (.A(_0180_),
    .B(_0184_),
    .X(_0187_));
 sky130_fd_sc_hd__nor2_1 _2186_ (.A(_0634_),
    .B(net65),
    .Y(_0188_));
 sky130_fd_sc_hd__and2b_1 _2187_ (.A_N(\pix_x[7] ),
    .B(\logo_left[7] ),
    .X(_0189_));
 sky130_fd_sc_hd__and2b_1 _2188_ (.A_N(\logo_left[7] ),
    .B(\pix_x[7] ),
    .X(_0190_));
 sky130_fd_sc_hd__inv_2 _2189_ (.A(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__or3_1 _2190_ (.A(_0188_),
    .B(_0189_),
    .C(_0190_),
    .X(_0192_));
 sky130_fd_sc_hd__nand2b_1 _2191_ (.A_N(\pix_x[8] ),
    .B(\logo_left[8] ),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2b_1 _2192_ (.A_N(\logo_left[8] ),
    .B(\pix_x[8] ),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _2193_ (.A(_0193_),
    .B(_0194_),
    .Y(_0195_));
 sky130_fd_sc_hd__a21oi_1 _2194_ (.A1(_0189_),
    .A2(_0195_),
    .B1(_0190_),
    .Y(_0196_));
 sky130_fd_sc_hd__o31a_1 _2195_ (.A1(_0634_),
    .A2(net63),
    .A3(_0196_),
    .B1(_0192_),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _2196_ (.A(_0519_),
    .B(net118),
    .X(_0198_));
 sky130_fd_sc_hd__xor2_1 _2197_ (.A(\logo_left[9] ),
    .B(\pix_x[9] ),
    .X(_0199_));
 sky130_fd_sc_hd__o22a_1 _2198_ (.A1(_0181_),
    .A2(_0198_),
    .B1(_0199_),
    .B2(_0193_),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _2199_ (.A1(_0181_),
    .A2(_0198_),
    .B1(_0199_),
    .B2(_0193_),
    .X(_0201_));
 sky130_fd_sc_hd__and4bb_1 _2200_ (.A_N(_0201_),
    .B_N(_0197_),
    .C(_0187_),
    .D(_0200_),
    .X(_0202_));
 sky130_fd_sc_hd__a21bo_1 _2201_ (.A1(_0191_),
    .A2(_0192_),
    .B1_N(_0195_),
    .X(_0203_));
 sky130_fd_sc_hd__o211a_1 _2202_ (.A1(_0183_),
    .A2(_0186_),
    .B1(_0202_),
    .C1(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__nor2_1 _2203_ (.A(net2),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__o21a_1 _2204_ (.A1(\pix_x[7] ),
    .A2(\pix_x[8] ),
    .B1(\pix_x[9] ),
    .X(_0206_));
 sky130_fd_sc_hd__or3_1 _2205_ (.A(_0532_),
    .B(\pix_y[9] ),
    .C(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__a211o_1 _2206_ (.A1(net118),
    .A2(_0536_),
    .B1(_0205_),
    .C1(_0207_),
    .X(_0208_));
 sky130_fd_sc_hd__o21ba_1 _2207_ (.A1(_1017_),
    .A2(_1140_),
    .B1_N(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__and2_1 _2208_ (.A(\logo_left[5] ),
    .B(net12),
    .X(_0210_));
 sky130_fd_sc_hd__nor2_1 _2209_ (.A(\logo_left[5] ),
    .B(net12),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_1 _2210_ (.A(_0210_),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__xnor2_1 _2211_ (.A(net52),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_1 _2212_ (.A(net130),
    .B(net41),
    .Y(_0214_));
 sky130_fd_sc_hd__xnor2_1 _2213_ (.A(\logo_left[4] ),
    .B(net42),
    .Y(_0215_));
 sky130_fd_sc_hd__o21a_1 _2214_ (.A1(net80),
    .A2(_0215_),
    .B1(_0214_),
    .X(_0216_));
 sky130_fd_sc_hd__xor2_1 _2215_ (.A(_0213_),
    .B(_0216_),
    .X(_0217_));
 sky130_fd_sc_hd__xnor2_1 _2216_ (.A(net80),
    .B(_0215_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_1 _2217_ (.A(\logo_left[3] ),
    .B(net88),
    .Y(_0219_));
 sky130_fd_sc_hd__or2_1 _2218_ (.A(\logo_left[3] ),
    .B(net88),
    .X(_0220_));
 sky130_fd_sc_hd__nand2_1 _2219_ (.A(_0219_),
    .B(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__o21a_1 _2220_ (.A1(_0676_),
    .A2(_0221_),
    .B1(_0219_),
    .X(_0222_));
 sky130_fd_sc_hd__nor2_1 _2221_ (.A(_0218_),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__xnor2_1 _2222_ (.A(net75),
    .B(_0221_),
    .Y(_0224_));
 sky130_fd_sc_hd__or2_1 _2223_ (.A(\logo_left[2] ),
    .B(_1018_),
    .X(_0225_));
 sky130_fd_sc_hd__and2b_1 _2224_ (.A_N(_0224_),
    .B(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__nand2_1 _2225_ (.A(\logo_left[2] ),
    .B(_1018_),
    .Y(_0227_));
 sky130_fd_sc_hd__a21oi_1 _2226_ (.A1(_0225_),
    .A2(_0227_),
    .B1(_0629_),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _2227_ (.A(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__xor2_1 _2228_ (.A(_0224_),
    .B(_0225_),
    .X(_0230_));
 sky130_fd_sc_hd__nor2_1 _2229_ (.A(_0229_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__and2_1 _2230_ (.A(_0218_),
    .B(_0222_),
    .X(_0232_));
 sky130_fd_sc_hd__nor2_1 _2231_ (.A(_0223_),
    .B(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__o21a_1 _2232_ (.A1(_0226_),
    .A2(_0231_),
    .B1(_0233_),
    .X(_0234_));
 sky130_fd_sc_hd__o21ai_1 _2233_ (.A1(_0223_),
    .A2(_0234_),
    .B1(_0217_),
    .Y(_0235_));
 sky130_fd_sc_hd__o21ai_1 _2234_ (.A1(_0213_),
    .A2(_0216_),
    .B1(_0235_),
    .Y(_0236_));
 sky130_fd_sc_hd__a21o_1 _2235_ (.A1(net52),
    .A2(_0212_),
    .B1(_0210_),
    .X(_0237_));
 sky130_fd_sc_hd__xnor2_1 _2236_ (.A(_0523_),
    .B(net27),
    .Y(_0238_));
 sky130_fd_sc_hd__xnor2_1 _2237_ (.A(net8),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__xnor2_1 _2238_ (.A(_0237_),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__xnor2_1 _2239_ (.A(_0236_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__mux2_1 _2240_ (.A0(\palette_inst.rrggbb[4] ),
    .A1(_0241_),
    .S(_0535_),
    .X(_0242_));
 sky130_fd_sc_hd__and3_1 _2241_ (.A(_0179_),
    .B(_0209_),
    .C(_0242_),
    .X(_0006_));
 sky130_fd_sc_hd__o211a_1 _2242_ (.A1(_0535_),
    .A2(net175),
    .B1(_0179_),
    .C1(_0209_),
    .X(_0007_));
 sky130_fd_sc_hd__nand2b_2 _2243_ (.A_N(\gamepad.driver.pmod_latch_prev ),
    .B(\gamepad.driver.pmod_latch_sync[1] ),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _2244_ (.A(net135),
    .B(net114),
    .Y(_0244_));
 sky130_fd_sc_hd__o22a_1 _2245_ (.A1(\gamepad.driver.shift_reg[0] ),
    .A2(net114),
    .B1(net104),
    .B2(net163),
    .X(_0008_));
 sky130_fd_sc_hd__o22a_1 _2246_ (.A1(\gamepad.driver.shift_reg[1] ),
    .A2(_0243_),
    .B1(net104),
    .B2(net167),
    .X(_0009_));
 sky130_fd_sc_hd__o22a_1 _2247_ (.A1(\gamepad.driver.shift_reg[2] ),
    .A2(_0243_),
    .B1(_0244_),
    .B2(net161),
    .X(_0010_));
 sky130_fd_sc_hd__o22a_1 _2248_ (.A1(\gamepad.driver.shift_reg[3] ),
    .A2(_0243_),
    .B1(_0244_),
    .B2(net173),
    .X(_0011_));
 sky130_fd_sc_hd__o22a_1 _2249_ (.A1(net183),
    .A2(net114),
    .B1(net104),
    .B2(net197),
    .X(_0012_));
 sky130_fd_sc_hd__o22a_1 _2250_ (.A1(net186),
    .A2(net114),
    .B1(net104),
    .B2(net194),
    .X(_0013_));
 sky130_fd_sc_hd__o22a_1 _2251_ (.A1(net188),
    .A2(net114),
    .B1(net104),
    .B2(net198),
    .X(_0014_));
 sky130_fd_sc_hd__o22a_1 _2252_ (.A1(net184),
    .A2(net114),
    .B1(net104),
    .B2(net207),
    .X(_0015_));
 sky130_fd_sc_hd__o22a_1 _2253_ (.A1(net180),
    .A2(net114),
    .B1(net104),
    .B2(net187),
    .X(_0016_));
 sky130_fd_sc_hd__o22a_1 _2254_ (.A1(\gamepad.driver.shift_reg[9] ),
    .A2(net114),
    .B1(net104),
    .B2(net165),
    .X(_0017_));
 sky130_fd_sc_hd__o22a_1 _2255_ (.A1(\gamepad.driver.shift_reg[10] ),
    .A2(net114),
    .B1(net104),
    .B2(net169),
    .X(_0018_));
 sky130_fd_sc_hd__o22a_1 _2256_ (.A1(\gamepad.driver.shift_reg[11] ),
    .A2(net114),
    .B1(net104),
    .B2(net159),
    .X(_0019_));
 sky130_fd_sc_hd__and4_1 _2257_ (.A(\gamepad.decoder.data_reg[9] ),
    .B(\gamepad.decoder.data_reg[8] ),
    .C(\gamepad.decoder.data_reg[11] ),
    .D(\gamepad.decoder.data_reg[10] ),
    .X(_0245_));
 sky130_fd_sc_hd__and4_1 _2258_ (.A(\gamepad.decoder.data_reg[5] ),
    .B(\gamepad.decoder.data_reg[4] ),
    .C(\gamepad.decoder.data_reg[7] ),
    .D(\gamepad.decoder.data_reg[6] ),
    .X(_0246_));
 sky130_fd_sc_hd__and4_1 _2259_ (.A(\gamepad.decoder.data_reg[1] ),
    .B(\gamepad.decoder.data_reg[0] ),
    .C(\gamepad.decoder.data_reg[3] ),
    .D(\gamepad.decoder.data_reg[2] ),
    .X(_0247_));
 sky130_fd_sc_hd__nand3_2 _2260_ (.A(_0245_),
    .B(_0246_),
    .C(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__and2_1 _2261_ (.A(\gamepad.decoder.data_reg[8] ),
    .B(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _2262_ (.A0(_0249_),
    .A1(gamepad_start_prev),
    .S(_0554_),
    .X(_0250_));
 sky130_fd_sc_hd__and2_1 _2263_ (.A(net133),
    .B(_0250_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _2264_ (.A(\pix_x[0] ),
    .B(\pix_x[1] ),
    .Y(_0251_));
 sky130_fd_sc_hd__nor2_1 _2265_ (.A(_0525_),
    .B(_0251_),
    .Y(_0252_));
 sky130_fd_sc_hd__and2_1 _2266_ (.A(\pix_x[3] ),
    .B(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__and3_1 _2267_ (.A(\pix_x[3] ),
    .B(\pix_x[4] ),
    .C(_0252_),
    .X(_0254_));
 sky130_fd_sc_hd__nand3b_1 _2268_ (.A_N(\pix_x[7] ),
    .B(\pix_x[8] ),
    .C(\pix_x[9] ),
    .Y(_0255_));
 sky130_fd_sc_hd__or4b_1 _2269_ (.A(\pix_x[5] ),
    .B(_0255_),
    .C(\pix_x[6] ),
    .D_N(_0254_),
    .X(_0256_));
 sky130_fd_sc_hd__inv_2 _2270_ (.A(_0256_),
    .Y(_0257_));
 sky130_fd_sc_hd__nor2_1 _2271_ (.A(_0532_),
    .B(_0257_),
    .Y(_0258_));
 sky130_fd_sc_hd__and2b_1 _2272_ (.A_N(net212),
    .B(net11),
    .X(_0021_));
 sky130_fd_sc_hd__or2_1 _2273_ (.A(\pix_x[0] ),
    .B(\pix_x[1] ),
    .X(_0259_));
 sky130_fd_sc_hd__and3_1 _2274_ (.A(_0251_),
    .B(net11),
    .C(_0259_),
    .X(_0022_));
 sky130_fd_sc_hd__a211oi_1 _2275_ (.A1(_0525_),
    .A2(_0251_),
    .B1(_0252_),
    .C1(_0532_),
    .Y(_0023_));
 sky130_fd_sc_hd__o21ai_1 _2276_ (.A1(\pix_x[3] ),
    .A2(_0252_),
    .B1(net134),
    .Y(_0260_));
 sky130_fd_sc_hd__nor2_1 _2277_ (.A(_0253_),
    .B(_0260_),
    .Y(_0024_));
 sky130_fd_sc_hd__o21ai_1 _2278_ (.A1(\pix_x[4] ),
    .A2(_0253_),
    .B1(net134),
    .Y(_0261_));
 sky130_fd_sc_hd__nor2_1 _2279_ (.A(_0254_),
    .B(_0261_),
    .Y(_0025_));
 sky130_fd_sc_hd__o21ai_1 _2280_ (.A1(\pix_x[5] ),
    .A2(_0254_),
    .B1(net11),
    .Y(_0262_));
 sky130_fd_sc_hd__a21oi_1 _2281_ (.A1(net213),
    .A2(_0254_),
    .B1(_0262_),
    .Y(_0026_));
 sky130_fd_sc_hd__a21o_1 _2282_ (.A1(\pix_x[5] ),
    .A2(_0254_),
    .B1(\pix_x[6] ),
    .X(_0263_));
 sky130_fd_sc_hd__and4_1 _2283_ (.A(\pix_x[4] ),
    .B(\pix_x[5] ),
    .C(\pix_x[6] ),
    .D(_0253_),
    .X(_0264_));
 sky130_fd_sc_hd__and3b_1 _2284_ (.A_N(_0264_),
    .B(net11),
    .C(_0263_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_1 _2285_ (.A(\pix_x[7] ),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__and2_1 _2286_ (.A(\pix_x[7] ),
    .B(_0264_),
    .X(_0266_));
 sky130_fd_sc_hd__and3b_1 _2287_ (.A_N(_0266_),
    .B(net10),
    .C(_0265_),
    .X(_0028_));
 sky130_fd_sc_hd__and3_1 _2288_ (.A(\pix_x[7] ),
    .B(\pix_x[8] ),
    .C(_0264_),
    .X(_0267_));
 sky130_fd_sc_hd__o21ai_1 _2289_ (.A1(\pix_x[8] ),
    .A2(_0266_),
    .B1(net11),
    .Y(_0268_));
 sky130_fd_sc_hd__nor2_1 _2290_ (.A(_0267_),
    .B(_0268_),
    .Y(_0029_));
 sky130_fd_sc_hd__o21ai_1 _2291_ (.A1(\pix_x[9] ),
    .A2(_0267_),
    .B1(net11),
    .Y(_0269_));
 sky130_fd_sc_hd__a21oi_1 _2292_ (.A1(net211),
    .A2(_0267_),
    .B1(_0269_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand2_1 _2293_ (.A(\gamepad.decoder.data_reg[5] ),
    .B(_0248_),
    .Y(_0270_));
 sky130_fd_sc_hd__or2_1 _2294_ (.A(\logo_left[1] ),
    .B(\logo_left[0] ),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _2295_ (.A(\logo_left[2] ),
    .B(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__or3_1 _2296_ (.A(\logo_left[7] ),
    .B(_0571_),
    .C(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__or2_1 _2297_ (.A(\logo_left[8] ),
    .B(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__o21bai_2 _2298_ (.A1(\logo_left[9] ),
    .A2(_0274_),
    .B1_N(_0270_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_1 _2299_ (.A(\gamepad.decoder.data_reg[4] ),
    .B(_0248_),
    .Y(_0276_));
 sky130_fd_sc_hd__or2_1 _2300_ (.A(\logo_left[9] ),
    .B(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__nor2_1 _2301_ (.A(_0580_),
    .B(_0277_),
    .Y(_0278_));
 sky130_fd_sc_hd__or2_2 _2302_ (.A(_0580_),
    .B(_0277_),
    .X(_0279_));
 sky130_fd_sc_hd__a31oi_4 _2303_ (.A1(net122),
    .A2(_0275_),
    .A3(_0279_),
    .B1(_0554_),
    .Y(_0280_));
 sky130_fd_sc_hd__a31o_2 _2304_ (.A1(net122),
    .A2(_0275_),
    .A3(_0279_),
    .B1(_0554_),
    .X(_0281_));
 sky130_fd_sc_hd__o21ai_1 _2305_ (.A1(\logo_left[0] ),
    .A2(_0280_),
    .B1(net135),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _2306_ (.A1(net210),
    .A2(_0280_),
    .B1(_0282_),
    .Y(_0031_));
 sky130_fd_sc_hd__a21o_1 _2307_ (.A1(_0576_),
    .A2(_0271_),
    .B1(_0279_),
    .X(_0283_));
 sky130_fd_sc_hd__nand2_1 _2308_ (.A(net123),
    .B(_0283_),
    .Y(_0284_));
 sky130_fd_sc_hd__a31o_1 _2309_ (.A1(_0576_),
    .A2(_0271_),
    .A3(_0279_),
    .B1(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _2310_ (.A(net115),
    .B(\logo_left[1] ),
    .X(_0286_));
 sky130_fd_sc_hd__and2_1 _2311_ (.A(net115),
    .B(\logo_left[1] ),
    .X(_0287_));
 sky130_fd_sc_hd__nand2_1 _2312_ (.A(net115),
    .B(\logo_left[1] ),
    .Y(_0288_));
 sky130_fd_sc_hd__and3_1 _2313_ (.A(\logo_left[0] ),
    .B(_0286_),
    .C(_0288_),
    .X(_0289_));
 sky130_fd_sc_hd__a21oi_1 _2314_ (.A1(_0286_),
    .A2(_0288_),
    .B1(\logo_left[0] ),
    .Y(_0290_));
 sky130_fd_sc_hd__o311a_1 _2315_ (.A1(net123),
    .A2(_0289_),
    .A3(_0290_),
    .B1(_0280_),
    .C1(_0285_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _2316_ (.A(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__o211a_1 _2317_ (.A1(\logo_left[1] ),
    .A2(_0280_),
    .B1(_0292_),
    .C1(net135),
    .X(_0032_));
 sky130_fd_sc_hd__nand2_1 _2318_ (.A(\logo_left[2] ),
    .B(_0271_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _2319_ (.A(_0272_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__xnor2_1 _2320_ (.A(_0283_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__xnor2_1 _2321_ (.A(dir_x),
    .B(\logo_left[2] ),
    .Y(_0296_));
 sky130_fd_sc_hd__o21a_1 _2322_ (.A1(_0287_),
    .A2(_0289_),
    .B1(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__nor3_1 _2323_ (.A(_0287_),
    .B(_0289_),
    .C(_0296_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _2324_ (.A(_0297_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand2_1 _2325_ (.A(_0524_),
    .B(_0281_),
    .Y(_0300_));
 sky130_fd_sc_hd__mux2_1 _2326_ (.A0(_0295_),
    .A1(_0299_),
    .S(net117),
    .X(_0301_));
 sky130_fd_sc_hd__o211a_1 _2327_ (.A1(_0281_),
    .A2(_0301_),
    .B1(_0300_),
    .C1(net135),
    .X(_0033_));
 sky130_fd_sc_hd__nand2_1 _2328_ (.A(net115),
    .B(\logo_left[3] ),
    .Y(_0302_));
 sky130_fd_sc_hd__or2_1 _2329_ (.A(_0518_),
    .B(\logo_left[3] ),
    .X(_0303_));
 sky130_fd_sc_hd__a21o_1 _2330_ (.A1(_0518_),
    .A2(\logo_left[2] ),
    .B1(_0297_),
    .X(_0304_));
 sky130_fd_sc_hd__a21oi_1 _2331_ (.A1(_0302_),
    .A2(_0303_),
    .B1(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__a31o_1 _2332_ (.A1(_0302_),
    .A2(_0303_),
    .A3(_0304_),
    .B1(net123),
    .X(_0306_));
 sky130_fd_sc_hd__and2_1 _2333_ (.A(_0577_),
    .B(_0278_),
    .X(_0307_));
 sky130_fd_sc_hd__o21bai_1 _2334_ (.A1(_0272_),
    .A2(_0278_),
    .B1_N(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nor2_1 _2335_ (.A(net131),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__a21o_1 _2336_ (.A1(net131),
    .A2(_0308_),
    .B1(net117),
    .X(_0310_));
 sky130_fd_sc_hd__o22a_1 _2337_ (.A1(_0305_),
    .A2(_0306_),
    .B1(_0309_),
    .B2(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__nor2_1 _2338_ (.A(_0281_),
    .B(_0311_),
    .Y(_0312_));
 sky130_fd_sc_hd__a211o_1 _2339_ (.A1(net131),
    .A2(_0281_),
    .B1(_0312_),
    .C1(_0532_),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_1 _2340_ (.A(_0518_),
    .B(net130),
    .Y(_0313_));
 sky130_fd_sc_hd__or2_1 _2341_ (.A(_0518_),
    .B(net130),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _2342_ (.A(_0313_),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_1 _2343_ (.A(_0303_),
    .B(_0304_),
    .Y(_0316_));
 sky130_fd_sc_hd__a21o_1 _2344_ (.A1(_0302_),
    .A2(_0316_),
    .B1(_0315_),
    .X(_0317_));
 sky130_fd_sc_hd__nand3_1 _2345_ (.A(_0302_),
    .B(_0315_),
    .C(_0316_),
    .Y(_0318_));
 sky130_fd_sc_hd__nand2_1 _2346_ (.A(_0317_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__or3_1 _2347_ (.A(net131),
    .B(_0272_),
    .C(_0278_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_1 _2348_ (.A(net131),
    .B(_0307_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21oi_1 _2349_ (.A1(_0320_),
    .A2(_0321_),
    .B1(net130),
    .Y(_0322_));
 sky130_fd_sc_hd__a31o_1 _2350_ (.A1(net130),
    .A2(_0320_),
    .A3(_0321_),
    .B1(net117),
    .X(_0323_));
 sky130_fd_sc_hd__a2bb2o_1 _2351_ (.A1_N(_0322_),
    .A2_N(_0323_),
    .B1(_0516_),
    .B2(_0319_),
    .X(_0324_));
 sky130_fd_sc_hd__nand2_1 _2352_ (.A(_0280_),
    .B(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__o211a_1 _2353_ (.A1(\logo_left[4] ),
    .A2(_0280_),
    .B1(_0325_),
    .C1(net135),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(_0320_),
    .A1(_0321_),
    .S(net130),
    .X(_0326_));
 sky130_fd_sc_hd__xnor2_1 _2355_ (.A(\logo_left[5] ),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__xor2_1 _2356_ (.A(dir_x),
    .B(\logo_left[5] ),
    .X(_0328_));
 sky130_fd_sc_hd__a21o_1 _2357_ (.A1(_0313_),
    .A2(_0317_),
    .B1(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__a31oi_1 _2358_ (.A1(_0313_),
    .A2(_0317_),
    .A3(_0328_),
    .B1(net123),
    .Y(_0330_));
 sky130_fd_sc_hd__a221o_1 _2359_ (.A1(net123),
    .A2(_0327_),
    .B1(_0329_),
    .B2(_0330_),
    .C1(_0281_),
    .X(_0331_));
 sky130_fd_sc_hd__o211a_1 _2360_ (.A1(\logo_left[5] ),
    .A2(_0280_),
    .B1(_0331_),
    .C1(net135),
    .X(_0036_));
 sky130_fd_sc_hd__xor2_1 _2361_ (.A(dir_x),
    .B(\logo_left[6] ),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _2362_ (.A(_0317_),
    .B(_0328_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _2363_ (.A(net115),
    .B(_0570_),
    .Y(_0334_));
 sky130_fd_sc_hd__and3_1 _2364_ (.A(_0332_),
    .B(_0333_),
    .C(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__a21oi_1 _2365_ (.A1(_0333_),
    .A2(_0334_),
    .B1(_0332_),
    .Y(_0336_));
 sky130_fd_sc_hd__or3_1 _2366_ (.A(net122),
    .B(_0335_),
    .C(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__o2bb2a_1 _2367_ (.A1_N(_0578_),
    .A2_N(_0307_),
    .B1(_0320_),
    .B2(_0570_),
    .X(_0338_));
 sky130_fd_sc_hd__o21ai_1 _2368_ (.A1(_0523_),
    .A2(_0338_),
    .B1(net123),
    .Y(_0339_));
 sky130_fd_sc_hd__a21o_1 _2369_ (.A1(_0523_),
    .A2(_0338_),
    .B1(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__a21oi_1 _2370_ (.A1(_0337_),
    .A2(_0340_),
    .B1(_0281_),
    .Y(_0341_));
 sky130_fd_sc_hd__a211o_1 _2371_ (.A1(\logo_left[6] ),
    .A2(_0281_),
    .B1(_0341_),
    .C1(_0532_),
    .X(_0037_));
 sky130_fd_sc_hd__xor2_1 _2372_ (.A(dir_x),
    .B(\logo_left[7] ),
    .X(_0342_));
 sky130_fd_sc_hd__a21oi_1 _2373_ (.A1(net115),
    .A2(\logo_left[6] ),
    .B1(_0336_),
    .Y(_0343_));
 sky130_fd_sc_hd__o21a_1 _2374_ (.A1(_0342_),
    .A2(_0343_),
    .B1(_0516_),
    .X(_0344_));
 sky130_fd_sc_hd__a21boi_1 _2375_ (.A1(_0342_),
    .A2(_0343_),
    .B1_N(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__nor2_1 _2376_ (.A(_0579_),
    .B(_0277_),
    .Y(_0346_));
 sky130_fd_sc_hd__a31o_1 _2377_ (.A1(\logo_left[6] ),
    .A2(_0577_),
    .A3(_0578_),
    .B1(\logo_left[7] ),
    .X(_0347_));
 sky130_fd_sc_hd__and3_1 _2378_ (.A(net122),
    .B(_0346_),
    .C(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_1 _2379_ (.A1(_0571_),
    .A2(_0272_),
    .B1(\logo_left[7] ),
    .Y(_0349_));
 sky130_fd_sc_hd__nand2_1 _2380_ (.A(_0273_),
    .B(_0349_),
    .Y(_0350_));
 sky130_fd_sc_hd__a31o_1 _2381_ (.A1(net122),
    .A2(_0279_),
    .A3(_0350_),
    .B1(_0348_),
    .X(_0351_));
 sky130_fd_sc_hd__o21a_1 _2382_ (.A1(_0345_),
    .A2(_0351_),
    .B1(_0280_),
    .X(_0352_));
 sky130_fd_sc_hd__a211o_1 _2383_ (.A1(\logo_left[7] ),
    .A2(_0281_),
    .B1(_0352_),
    .C1(_0532_),
    .X(_0038_));
 sky130_fd_sc_hd__or2_1 _2384_ (.A(net115),
    .B(\logo_left[8] ),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_1 _2385_ (.A(net115),
    .B(\logo_left[8] ),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _2386_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__or3_1 _2387_ (.A(_0332_),
    .B(_0333_),
    .C(_0342_),
    .X(_0356_));
 sky130_fd_sc_hd__o21ai_1 _2388_ (.A1(\logo_left[7] ),
    .A2(\logo_left[6] ),
    .B1(net115),
    .Y(_0357_));
 sky130_fd_sc_hd__and3_1 _2389_ (.A(_0334_),
    .B(_0356_),
    .C(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__a21o_1 _2390_ (.A1(_0355_),
    .A2(_0358_),
    .B1(net122),
    .X(_0359_));
 sky130_fd_sc_hd__o21ba_1 _2391_ (.A1(_0355_),
    .A2(_0358_),
    .B1_N(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__a21o_1 _2392_ (.A1(_0273_),
    .A2(_0279_),
    .B1(_0346_),
    .X(_0361_));
 sky130_fd_sc_hd__xnor2_1 _2393_ (.A(\logo_left[8] ),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__a21o_1 _2394_ (.A1(net122),
    .A2(_0362_),
    .B1(_0281_),
    .X(_0363_));
 sky130_fd_sc_hd__o221a_1 _2395_ (.A1(\logo_left[8] ),
    .A2(_0280_),
    .B1(_0360_),
    .B2(_0363_),
    .C1(net134),
    .X(_0039_));
 sky130_fd_sc_hd__o21ai_1 _2396_ (.A1(_0355_),
    .A2(_0358_),
    .B1(_0354_),
    .Y(_0364_));
 sky130_fd_sc_hd__nand2_1 _2397_ (.A(dir_x),
    .B(\logo_left[9] ),
    .Y(_0365_));
 sky130_fd_sc_hd__nand2_1 _2398_ (.A(_0573_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__xnor2_1 _2399_ (.A(_0364_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__nor2_1 _2400_ (.A(net122),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__xnor2_1 _2401_ (.A(\logo_left[9] ),
    .B(_0274_),
    .Y(_0369_));
 sky130_fd_sc_hd__a31o_1 _2402_ (.A1(net122),
    .A2(_0279_),
    .A3(_0369_),
    .B1(_0281_),
    .X(_0370_));
 sky130_fd_sc_hd__o221a_1 _2403_ (.A1(\logo_left[9] ),
    .A2(_0280_),
    .B1(_0368_),
    .B2(_0370_),
    .C1(net134),
    .X(_0040_));
 sky130_fd_sc_hd__nand2_1 _2404_ (.A(\gamepad.decoder.data_reg[7] ),
    .B(_0248_),
    .Y(_0371_));
 sky130_fd_sc_hd__or2_2 _2405_ (.A(\logo_top[1] ),
    .B(\logo_top[0] ),
    .X(_0372_));
 sky130_fd_sc_hd__inv_2 _2406_ (.A(_0372_),
    .Y(_0373_));
 sky130_fd_sc_hd__or4b_2 _2407_ (.A(\logo_top[8] ),
    .B(_0372_),
    .C(net125),
    .D_N(_0568_),
    .X(_0374_));
 sky130_fd_sc_hd__inv_2 _2408_ (.A(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__o21bai_2 _2409_ (.A1(\logo_top[9] ),
    .A2(_0374_),
    .B1_N(_0371_),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _2410_ (.A(\gamepad.decoder.data_reg[6] ),
    .B(_0248_),
    .Y(_0377_));
 sky130_fd_sc_hd__a21o_1 _2411_ (.A1(\logo_top[6] ),
    .A2(\logo_top[5] ),
    .B1(net125),
    .X(_0378_));
 sky130_fd_sc_hd__a211o_1 _2412_ (.A1(\logo_top[8] ),
    .A2(_0378_),
    .B1(_0377_),
    .C1(\logo_top[9] ),
    .X(_0379_));
 sky130_fd_sc_hd__nor2_1 _2413_ (.A(_0563_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__or2_2 _2414_ (.A(_0563_),
    .B(_0379_),
    .X(_0381_));
 sky130_fd_sc_hd__a31oi_4 _2415_ (.A1(net121),
    .A2(_0376_),
    .A3(_0381_),
    .B1(_0554_),
    .Y(_0382_));
 sky130_fd_sc_hd__a31o_1 _2416_ (.A1(net121),
    .A2(_0376_),
    .A3(_0381_),
    .B1(_0554_),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _2417_ (.A1(\logo_top[0] ),
    .A2(_0382_),
    .B1(_0532_),
    .Y(_0384_));
 sky130_fd_sc_hd__o21a_1 _2418_ (.A1(\logo_top[0] ),
    .A2(_0382_),
    .B1(_0384_),
    .X(_0041_));
 sky130_fd_sc_hd__a21o_1 _2419_ (.A1(_0556_),
    .A2(_0372_),
    .B1(_0381_),
    .X(_0385_));
 sky130_fd_sc_hd__nand3_1 _2420_ (.A(_0556_),
    .B(_0372_),
    .C(_0381_),
    .Y(_0386_));
 sky130_fd_sc_hd__or2_1 _2421_ (.A(net116),
    .B(\logo_top[1] ),
    .X(_0387_));
 sky130_fd_sc_hd__and2_1 _2422_ (.A(net116),
    .B(\logo_top[1] ),
    .X(_0388_));
 sky130_fd_sc_hd__nand2_1 _2423_ (.A(net116),
    .B(\logo_top[1] ),
    .Y(_0389_));
 sky130_fd_sc_hd__and3_1 _2424_ (.A(\logo_top[0] ),
    .B(_0387_),
    .C(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__a21oi_1 _2425_ (.A1(_0387_),
    .A2(_0389_),
    .B1(\logo_top[0] ),
    .Y(_0391_));
 sky130_fd_sc_hd__nor3_1 _2426_ (.A(net121),
    .B(_0390_),
    .C(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__a311o_1 _2427_ (.A1(net120),
    .A2(_0385_),
    .A3(_0386_),
    .B1(_0392_),
    .C1(_0383_),
    .X(_0393_));
 sky130_fd_sc_hd__o211a_1 _2428_ (.A1(\logo_top[1] ),
    .A2(_0382_),
    .B1(_0393_),
    .C1(net133),
    .X(_0042_));
 sky130_fd_sc_hd__xor2_1 _2429_ (.A(\logo_top[2] ),
    .B(_0372_),
    .X(_0394_));
 sky130_fd_sc_hd__xnor2_1 _2430_ (.A(_0385_),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__xnor2_1 _2431_ (.A(net124),
    .B(\logo_top[2] ),
    .Y(_0396_));
 sky130_fd_sc_hd__nor3_1 _2432_ (.A(_0388_),
    .B(_0390_),
    .C(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__o21a_1 _2433_ (.A1(_0388_),
    .A2(_0390_),
    .B1(_0396_),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _2434_ (.A(\logo_top[2] ),
    .B(_0382_),
    .X(_0399_));
 sky130_fd_sc_hd__nor3_1 _2435_ (.A(net120),
    .B(_0397_),
    .C(_0398_),
    .Y(_0400_));
 sky130_fd_sc_hd__nor2_1 _2436_ (.A(net117),
    .B(_0395_),
    .Y(_0401_));
 sky130_fd_sc_hd__o311a_1 _2437_ (.A1(net9),
    .A2(_0400_),
    .A3(_0401_),
    .B1(_0399_),
    .C1(net133),
    .X(_0043_));
 sky130_fd_sc_hd__or2_1 _2438_ (.A(net116),
    .B(net129),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _2439_ (.A(_0517_),
    .B(net129),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _2440_ (.A(_0402_),
    .B(_0403_),
    .Y(_0404_));
 sky130_fd_sc_hd__a21oi_1 _2441_ (.A1(net116),
    .A2(\logo_top[2] ),
    .B1(_0398_),
    .Y(_0405_));
 sky130_fd_sc_hd__xnor2_1 _2442_ (.A(_0404_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__or3_1 _2443_ (.A(\logo_top[2] ),
    .B(_0372_),
    .C(_0380_),
    .X(_0407_));
 sky130_fd_sc_hd__a21bo_1 _2444_ (.A1(_0557_),
    .A2(_0380_),
    .B1_N(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__nor2_1 _2445_ (.A(net129),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__a21o_1 _2446_ (.A1(net129),
    .A2(_0408_),
    .B1(net117),
    .X(_0410_));
 sky130_fd_sc_hd__o22a_1 _2447_ (.A1(net120),
    .A2(_0406_),
    .B1(_0409_),
    .B2(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__nor2_1 _2448_ (.A(net9),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__a211o_1 _2449_ (.A1(net129),
    .A2(net9),
    .B1(_0412_),
    .C1(_0532_),
    .X(_0044_));
 sky130_fd_sc_hd__and3_1 _2450_ (.A(net129),
    .B(_0557_),
    .C(_0380_),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _2451_ (.A(\logo_top[3] ),
    .B(_0407_),
    .Y(_0414_));
 sky130_fd_sc_hd__or3_1 _2452_ (.A(net128),
    .B(_0413_),
    .C(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__o21ai_1 _2453_ (.A1(_0413_),
    .A2(_0414_),
    .B1(net128),
    .Y(_0416_));
 sky130_fd_sc_hd__and3_1 _2454_ (.A(net120),
    .B(_0415_),
    .C(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _2455_ (.A(net116),
    .B(net128),
    .Y(_0418_));
 sky130_fd_sc_hd__or2_1 _2456_ (.A(net116),
    .B(net128),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _2457_ (.A1(_0517_),
    .A2(_0565_),
    .B1(_0398_),
    .B2(_0402_),
    .X(_0420_));
 sky130_fd_sc_hd__a21o_1 _2458_ (.A1(_0418_),
    .A2(_0419_),
    .B1(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__nand3_1 _2459_ (.A(_0418_),
    .B(_0419_),
    .C(_0420_),
    .Y(_0422_));
 sky130_fd_sc_hd__a31o_1 _2460_ (.A1(net117),
    .A2(_0421_),
    .A3(_0422_),
    .B1(net9),
    .X(_0423_));
 sky130_fd_sc_hd__o221a_1 _2461_ (.A1(net128),
    .A2(_0382_),
    .B1(_0417_),
    .B2(_0423_),
    .C1(net133),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _2462_ (.A(_0558_),
    .B(_0380_),
    .X(_0424_));
 sky130_fd_sc_hd__and2b_1 _2463_ (.A_N(net128),
    .B(_0414_),
    .X(_0425_));
 sky130_fd_sc_hd__o21ai_1 _2464_ (.A1(_0424_),
    .A2(_0425_),
    .B1(net127),
    .Y(_0426_));
 sky130_fd_sc_hd__o31a_1 _2465_ (.A1(net127),
    .A2(_0424_),
    .A3(_0425_),
    .B1(net120),
    .X(_0427_));
 sky130_fd_sc_hd__nand2_1 _2466_ (.A(_0418_),
    .B(_0422_),
    .Y(_0428_));
 sky130_fd_sc_hd__xor2_1 _2467_ (.A(net124),
    .B(net127),
    .X(_0429_));
 sky130_fd_sc_hd__xnor2_1 _2468_ (.A(_0428_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_1 _2469_ (.A(_0522_),
    .B(net9),
    .Y(_0431_));
 sky130_fd_sc_hd__a22o_1 _2470_ (.A1(_0426_),
    .A2(_0427_),
    .B1(_0430_),
    .B2(net117),
    .X(_0432_));
 sky130_fd_sc_hd__o211a_1 _2471_ (.A1(net9),
    .A2(_0432_),
    .B1(_0431_),
    .C1(net133),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_1 _2472_ (.A1(_0566_),
    .A2(_0414_),
    .B1(_0424_),
    .B2(net127),
    .X(_0433_));
 sky130_fd_sc_hd__a21oi_1 _2473_ (.A1(net126),
    .A2(_0433_),
    .B1(net117),
    .Y(_0434_));
 sky130_fd_sc_hd__o21a_1 _2474_ (.A1(net126),
    .A2(_0433_),
    .B1(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__xnor2_1 _2475_ (.A(net124),
    .B(net126),
    .Y(_0436_));
 sky130_fd_sc_hd__nor2_1 _2476_ (.A(_0422_),
    .B(_0429_),
    .Y(_0437_));
 sky130_fd_sc_hd__nor2_1 _2477_ (.A(net124),
    .B(_0566_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor3_1 _2478_ (.A(_0436_),
    .B(_0437_),
    .C(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__o21a_1 _2479_ (.A1(_0437_),
    .A2(_0438_),
    .B1(_0436_),
    .X(_0440_));
 sky130_fd_sc_hd__o31ai_1 _2480_ (.A1(net120),
    .A2(_0439_),
    .A3(_0440_),
    .B1(_0382_),
    .Y(_0441_));
 sky130_fd_sc_hd__a2bb2o_1 _2481_ (.A1_N(_0435_),
    .A2_N(_0441_),
    .B1(_0521_),
    .B2(net9),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_1 _2482_ (.A(net133),
    .B(_0442_),
    .Y(_0047_));
 sky130_fd_sc_hd__xor2_1 _2483_ (.A(net124),
    .B(net125),
    .X(_0443_));
 sky130_fd_sc_hd__a21oi_1 _2484_ (.A1(net116),
    .A2(net126),
    .B1(_0440_),
    .Y(_0444_));
 sky130_fd_sc_hd__xnor2_1 _2485_ (.A(_0443_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__and3_1 _2486_ (.A(_0568_),
    .B(_0373_),
    .C(_0381_),
    .X(_0446_));
 sky130_fd_sc_hd__a31o_1 _2487_ (.A1(net126),
    .A2(net127),
    .A3(_0424_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _2488_ (.A(\logo_top[7] ),
    .B(_0447_),
    .Y(_0448_));
 sky130_fd_sc_hd__o21a_1 _2489_ (.A1(\logo_top[7] ),
    .A2(_0447_),
    .B1(net120),
    .X(_0449_));
 sky130_fd_sc_hd__o2bb2a_1 _2490_ (.A1_N(_0449_),
    .A2_N(_0448_),
    .B1(_0445_),
    .B2(net120),
    .X(_0450_));
 sky130_fd_sc_hd__nor2_1 _2491_ (.A(net9),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__a211o_1 _2492_ (.A1(net125),
    .A2(net9),
    .B1(_0451_),
    .C1(_0532_),
    .X(_0048_));
 sky130_fd_sc_hd__a21oi_1 _2493_ (.A1(_0520_),
    .A2(_0566_),
    .B1(net124),
    .Y(_0452_));
 sky130_fd_sc_hd__o211a_1 _2494_ (.A1(net116),
    .A2(\logo_top[7] ),
    .B1(_0436_),
    .C1(_0437_),
    .X(_0453_));
 sky130_fd_sc_hd__a211o_1 _2495_ (.A1(net116),
    .A2(net126),
    .B1(_0452_),
    .C1(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__nand2_1 _2496_ (.A(net124),
    .B(\logo_top[8] ),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_1 _2497_ (.A(_0569_),
    .B(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__nand2_1 _2498_ (.A(_0454_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__or2_1 _2499_ (.A(_0454_),
    .B(_0456_),
    .X(_0458_));
 sky130_fd_sc_hd__and3_1 _2500_ (.A(net117),
    .B(_0457_),
    .C(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__o41a_1 _2501_ (.A1(net125),
    .A2(\logo_top[6] ),
    .A3(_0567_),
    .A4(_0372_),
    .B1(\logo_top[8] ),
    .X(_0460_));
 sky130_fd_sc_hd__o32a_1 _2502_ (.A1(_0375_),
    .A2(_0380_),
    .A3(_0460_),
    .B1(_0379_),
    .B2(_0560_),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_1 _2503_ (.A1(net120),
    .A2(_0461_),
    .B1(net9),
    .X(_0462_));
 sky130_fd_sc_hd__o221a_1 _2504_ (.A1(\logo_top[8] ),
    .A2(_0382_),
    .B1(_0459_),
    .B2(_0462_),
    .C1(net133),
    .X(_0049_));
 sky130_fd_sc_hd__o211ai_1 _2505_ (.A1(_0438_),
    .A2(_0453_),
    .B1(net124),
    .C1(\logo_top[8] ),
    .Y(_0463_));
 sky130_fd_sc_hd__o21ai_1 _2506_ (.A1(_0569_),
    .A2(_0454_),
    .B1(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__a21oi_1 _2507_ (.A1(\logo_top[9] ),
    .A2(_0464_),
    .B1(net121),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_1 _2508_ (.A1(\logo_top[9] ),
    .A2(_0464_),
    .B1(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__xnor2_1 _2509_ (.A(\logo_top[9] ),
    .B(_0374_),
    .Y(_0467_));
 sky130_fd_sc_hd__a31o_1 _2510_ (.A1(net121),
    .A2(_0381_),
    .A3(_0467_),
    .B1(_0383_),
    .X(_0468_));
 sky130_fd_sc_hd__o221a_1 _2511_ (.A1(\logo_top[9] ),
    .A2(_0382_),
    .B1(_0466_),
    .B2(_0468_),
    .C1(net133),
    .X(_0050_));
 sky130_fd_sc_hd__a31o_1 _2512_ (.A1(_0585_),
    .A2(_0270_),
    .A3(_0276_),
    .B1(_0555_),
    .X(_0469_));
 sky130_fd_sc_hd__nand2b_1 _2513_ (.A_N(_0270_),
    .B(_0575_),
    .Y(_0470_));
 sky130_fd_sc_hd__o21ai_1 _2514_ (.A1(\logo_left[9] ),
    .A2(_0584_),
    .B1(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__mux2_1 _2515_ (.A0(_0471_),
    .A1(net115),
    .S(_0469_),
    .X(_0472_));
 sky130_fd_sc_hd__nand2_1 _2516_ (.A(net134),
    .B(_0472_),
    .Y(_0051_));
 sky130_fd_sc_hd__and3_1 _2517_ (.A(_0564_),
    .B(_0587_),
    .C(_0371_),
    .X(_0473_));
 sky130_fd_sc_hd__a21oi_1 _2518_ (.A1(_0377_),
    .A2(_0473_),
    .B1(_0555_),
    .Y(_0474_));
 sky130_fd_sc_hd__a32o_1 _2519_ (.A1(\gamepad.decoder.data_reg[7] ),
    .A2(_0587_),
    .A3(_0248_),
    .B1(_0563_),
    .B2(dir_y),
    .X(_0475_));
 sky130_fd_sc_hd__nand2_1 _2520_ (.A(_0474_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__o211a_1 _2521_ (.A1(net124),
    .A2(_0474_),
    .B1(_0476_),
    .C1(net133),
    .X(_0052_));
 sky130_fd_sc_hd__or3b_1 _2522_ (.A(gamepad_start_prev),
    .B(_0554_),
    .C_N(_0249_),
    .X(_0477_));
 sky130_fd_sc_hd__xnor2_1 _2523_ (.A(net117),
    .B(_0477_),
    .Y(_0478_));
 sky130_fd_sc_hd__nor2_1 _2524_ (.A(_0532_),
    .B(_0478_),
    .Y(_0053_));
 sky130_fd_sc_hd__mux2_1 _2525_ (.A0(net202),
    .A1(\pix_y[0] ),
    .S(net132),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _2526_ (.A0(net209),
    .A1(net119),
    .S(net132),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _2527_ (.A0(net205),
    .A1(\pix_y[2] ),
    .S(net132),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _2528_ (.A0(net203),
    .A1(\pix_y[3] ),
    .S(net132),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _2529_ (.A0(net196),
    .A1(\pix_y[4] ),
    .S(net132),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _2530_ (.A0(net193),
    .A1(\pix_y[5] ),
    .S(net132),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _2531_ (.A0(net200),
    .A1(\pix_y[6] ),
    .S(net132),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _2532_ (.A0(net204),
    .A1(\pix_y[7] ),
    .S(net132),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _2533_ (.A0(net201),
    .A1(net118),
    .S(net132),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _2534_ (.A0(net195),
    .A1(\pix_y[9] ),
    .S(net132),
    .X(_0066_));
 sky130_fd_sc_hd__and3_1 _2535_ (.A(net99),
    .B(_0225_),
    .C(_0227_),
    .X(_0479_));
 sky130_fd_sc_hd__nor2_1 _2536_ (.A(_0228_),
    .B(_0479_),
    .Y(_0480_));
 sky130_fd_sc_hd__mux2_1 _2537_ (.A0(\palette_inst.rrggbb[0] ),
    .A1(_0480_),
    .S(_0535_),
    .X(_0481_));
 sky130_fd_sc_hd__and3_1 _2538_ (.A(_0179_),
    .B(_0209_),
    .C(_0481_),
    .X(_0067_));
 sky130_fd_sc_hd__and2_1 _2539_ (.A(_0229_),
    .B(_0230_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_1 _2540_ (.A(_0231_),
    .B(_0482_),
    .Y(_0483_));
 sky130_fd_sc_hd__mux2_1 _2541_ (.A0(\palette_inst.rrggbb[1] ),
    .A1(_0483_),
    .S(_0535_),
    .X(_0484_));
 sky130_fd_sc_hd__and3_1 _2542_ (.A(_0179_),
    .B(_0209_),
    .C(_0484_),
    .X(_0068_));
 sky130_fd_sc_hd__or3_1 _2543_ (.A(_0226_),
    .B(_0231_),
    .C(_0233_),
    .X(_0485_));
 sky130_fd_sc_hd__nor2_1 _2544_ (.A(net3),
    .B(_0234_),
    .Y(_0486_));
 sky130_fd_sc_hd__a22o_1 _2545_ (.A1(net3),
    .A2(\palette_inst.rrggbb[2] ),
    .B1(_0485_),
    .B2(_0486_),
    .X(_0487_));
 sky130_fd_sc_hd__and3_1 _2546_ (.A(_0179_),
    .B(_0209_),
    .C(_0487_),
    .X(_0069_));
 sky130_fd_sc_hd__or3_1 _2547_ (.A(_0217_),
    .B(_0223_),
    .C(_0234_),
    .X(_0488_));
 sky130_fd_sc_hd__a21o_1 _2548_ (.A1(_0235_),
    .A2(_0488_),
    .B1(net3),
    .X(_0489_));
 sky130_fd_sc_hd__o2111a_1 _2549_ (.A1(_0535_),
    .A2(net182),
    .B1(_0179_),
    .C1(_0209_),
    .D1(_0489_),
    .X(_0070_));
 sky130_fd_sc_hd__nand2b_1 _2550_ (.A_N(\gamepad.driver.pmod_clk_prev ),
    .B(\gamepad.driver.pmod_clk_sync[1] ),
    .Y(_0490_));
 sky130_fd_sc_hd__nand2_1 _2551_ (.A(net135),
    .B(_0490_),
    .Y(_0491_));
 sky130_fd_sc_hd__o22a_1 _2552_ (.A1(net171),
    .A2(_0490_),
    .B1(_0491_),
    .B2(\gamepad.driver.shift_reg[0] ),
    .X(_0071_));
 sky130_fd_sc_hd__o22a_1 _2553_ (.A1(\gamepad.driver.shift_reg[0] ),
    .A2(_0490_),
    .B1(_0491_),
    .B2(net191),
    .X(_0072_));
 sky130_fd_sc_hd__o22a_1 _2554_ (.A1(net191),
    .A2(net113),
    .B1(net103),
    .B2(net199),
    .X(_0073_));
 sky130_fd_sc_hd__o22a_1 _2555_ (.A1(\gamepad.driver.shift_reg[2] ),
    .A2(net113),
    .B1(net103),
    .B2(net178),
    .X(_0074_));
 sky130_fd_sc_hd__o22a_1 _2556_ (.A1(net178),
    .A2(net113),
    .B1(net103),
    .B2(net183),
    .X(_0075_));
 sky130_fd_sc_hd__o22a_1 _2557_ (.A1(net183),
    .A2(net113),
    .B1(net103),
    .B2(net186),
    .X(_0076_));
 sky130_fd_sc_hd__o22a_1 _2558_ (.A1(net186),
    .A2(net113),
    .B1(net103),
    .B2(net188),
    .X(_0077_));
 sky130_fd_sc_hd__o22a_1 _2559_ (.A1(\gamepad.driver.shift_reg[6] ),
    .A2(net113),
    .B1(net103),
    .B2(net184),
    .X(_0078_));
 sky130_fd_sc_hd__o22a_1 _2560_ (.A1(\gamepad.driver.shift_reg[7] ),
    .A2(net113),
    .B1(net103),
    .B2(net180),
    .X(_0079_));
 sky130_fd_sc_hd__o22a_1 _2561_ (.A1(net180),
    .A2(net113),
    .B1(net103),
    .B2(net189),
    .X(_0080_));
 sky130_fd_sc_hd__o22a_1 _2562_ (.A1(net189),
    .A2(net113),
    .B1(net103),
    .B2(net190),
    .X(_0081_));
 sky130_fd_sc_hd__o22a_1 _2563_ (.A1(\gamepad.driver.shift_reg[10] ),
    .A2(net113),
    .B1(net103),
    .B2(net176),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _2564_ (.A(net136),
    .B(net6),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _2565_ (.A(net136),
    .B(net157),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _2566_ (.A(net136),
    .B(net5),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _2567_ (.A(net136),
    .B(net158),
    .X(_0086_));
 sky130_fd_sc_hd__and2_1 _2568_ (.A(net136),
    .B(net4),
    .X(_0087_));
 sky130_fd_sc_hd__and2_1 _2569_ (.A(net136),
    .B(net156),
    .X(_0088_));
 sky130_fd_sc_hd__or4_1 _2570_ (.A(\pix_y[0] ),
    .B(\pix_y[1] ),
    .C(_0528_),
    .D(net118),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _2571_ (.A(\pix_y[3] ),
    .B(\pix_y[9] ),
    .Y(_0493_));
 sky130_fd_sc_hd__o311a_2 _2572_ (.A1(_0551_),
    .A2(_0492_),
    .A3(_0493_),
    .B1(_0257_),
    .C1(net137),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _2573_ (.A0(net10),
    .A1(_0494_),
    .S(_0526_),
    .X(_0089_));
 sky130_fd_sc_hd__xor2_1 _2574_ (.A(\pix_y[0] ),
    .B(net119),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _2575_ (.A1(net119),
    .A2(net10),
    .B1(_0494_),
    .B2(_0495_),
    .X(_0090_));
 sky130_fd_sc_hd__a21oi_1 _2576_ (.A1(\pix_y[0] ),
    .A2(net119),
    .B1(\pix_y[2] ),
    .Y(_0496_));
 sky130_fd_sc_hd__and3_1 _2577_ (.A(\pix_y[0] ),
    .B(net119),
    .C(\pix_y[2] ),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_1 _2578_ (.A(_0496_),
    .B(_0497_),
    .Y(_0498_));
 sky130_fd_sc_hd__a22o_1 _2579_ (.A1(\pix_y[2] ),
    .A2(net10),
    .B1(_0494_),
    .B2(_0498_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _2580_ (.A(\pix_y[3] ),
    .B(_0497_),
    .Y(_0499_));
 sky130_fd_sc_hd__and2_1 _2581_ (.A(\pix_y[3] ),
    .B(_0497_),
    .X(_0500_));
 sky130_fd_sc_hd__nor2_1 _2582_ (.A(_0499_),
    .B(_0500_),
    .Y(_0501_));
 sky130_fd_sc_hd__a22o_1 _2583_ (.A1(net214),
    .A2(net10),
    .B1(_0494_),
    .B2(_0501_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_1 _2584_ (.A(\pix_y[4] ),
    .B(_0500_),
    .Y(_0502_));
 sky130_fd_sc_hd__and3_1 _2585_ (.A(\pix_y[3] ),
    .B(\pix_y[4] ),
    .C(_0497_),
    .X(_0503_));
 sky130_fd_sc_hd__nor2_1 _2586_ (.A(_0502_),
    .B(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__a22o_1 _2587_ (.A1(\pix_y[4] ),
    .A2(net10),
    .B1(_0494_),
    .B2(_0504_),
    .X(_0093_));
 sky130_fd_sc_hd__xnor2_1 _2588_ (.A(_0531_),
    .B(_0503_),
    .Y(_0505_));
 sky130_fd_sc_hd__a22o_1 _2589_ (.A1(\pix_y[5] ),
    .A2(net10),
    .B1(_0494_),
    .B2(_0505_),
    .X(_0094_));
 sky130_fd_sc_hd__a21oi_1 _2590_ (.A1(\pix_y[5] ),
    .A2(_0503_),
    .B1(\pix_y[6] ),
    .Y(_0506_));
 sky130_fd_sc_hd__and3_1 _2591_ (.A(\pix_y[5] ),
    .B(\pix_y[6] ),
    .C(_0503_),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_1 _2592_ (.A(_0506_),
    .B(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__a22o_1 _2593_ (.A1(\pix_y[6] ),
    .A2(net10),
    .B1(_0494_),
    .B2(_0508_),
    .X(_0095_));
 sky130_fd_sc_hd__or2_1 _2594_ (.A(\pix_y[7] ),
    .B(_0507_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2_1 _2595_ (.A(\pix_y[7] ),
    .B(_0507_),
    .Y(_0510_));
 sky130_fd_sc_hd__a32o_1 _2596_ (.A1(_0494_),
    .A2(_0509_),
    .A3(_0510_),
    .B1(net10),
    .B2(\pix_y[7] ),
    .X(_0096_));
 sky130_fd_sc_hd__nand3_1 _2597_ (.A(net118),
    .B(\pix_y[7] ),
    .C(_0507_),
    .Y(_0511_));
 sky130_fd_sc_hd__a21o_1 _2598_ (.A1(_0494_),
    .A2(_0511_),
    .B1(net10),
    .X(_0512_));
 sky130_fd_sc_hd__and3_1 _2599_ (.A(\pix_y[7] ),
    .B(_0494_),
    .C(_0507_),
    .X(_0513_));
 sky130_fd_sc_hd__o21a_1 _2600_ (.A1(net118),
    .A2(_0513_),
    .B1(_0512_),
    .X(_0097_));
 sky130_fd_sc_hd__and3b_1 _2601_ (.A_N(\pix_y[9] ),
    .B(_0513_),
    .C(net118),
    .X(_0514_));
 sky130_fd_sc_hd__a21o_1 _2602_ (.A1(\pix_y[9] ),
    .A2(_0512_),
    .B1(_0514_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _2603_ (.A(_0055_),
    .B(_0100_),
    .X(_0099_));
 sky130_fd_sc_hd__dfxtp_2 _2604_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0006_),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__dfxtp_2 _2605_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0007_),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__dfxtp_1 _2606_ (.CLK(clknet_3_4__leaf_clk),
    .D(net164),
    .Q(\gamepad.decoder.data_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2607_ (.CLK(clknet_3_4__leaf_clk),
    .D(net168),
    .Q(\gamepad.decoder.data_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2608_ (.CLK(clknet_3_4__leaf_clk),
    .D(net162),
    .Q(\gamepad.decoder.data_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2609_ (.CLK(clknet_3_7__leaf_clk),
    .D(net174),
    .Q(\gamepad.decoder.data_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2610_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0012_),
    .Q(\gamepad.decoder.data_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2611_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0013_),
    .Q(\gamepad.decoder.data_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2612_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0014_),
    .Q(\gamepad.decoder.data_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2613_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0015_),
    .Q(\gamepad.decoder.data_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2614_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0016_),
    .Q(\gamepad.decoder.data_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2615_ (.CLK(clknet_3_6__leaf_clk),
    .D(net166),
    .Q(\gamepad.decoder.data_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2616_ (.CLK(clknet_3_7__leaf_clk),
    .D(net170),
    .Q(\gamepad.decoder.data_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2617_ (.CLK(clknet_3_6__leaf_clk),
    .D(net160),
    .Q(\gamepad.decoder.data_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2618_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0020_),
    .Q(gamepad_start_prev));
 sky130_fd_sc_hd__dfxtp_1 _2619_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0021_),
    .Q(\pix_x[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2620_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0022_),
    .Q(\pix_x[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2621_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0023_),
    .Q(\pix_x[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2622_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0024_),
    .Q(\pix_x[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2623_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0025_),
    .Q(\pix_x[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2624_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0026_),
    .Q(\pix_x[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2625_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0027_),
    .Q(\pix_x[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2626_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0028_),
    .Q(\pix_x[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2627_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0029_),
    .Q(\pix_x[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2628_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0030_),
    .Q(\pix_x[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2629_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0031_),
    .Q(\logo_left[0] ));
 sky130_fd_sc_hd__dfxtp_2 _2630_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0032_),
    .Q(\logo_left[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2631_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0033_),
    .Q(\logo_left[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2632_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0034_),
    .Q(\logo_left[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2633_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0035_),
    .Q(\logo_left[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2634_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0036_),
    .Q(\logo_left[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2635_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0037_),
    .Q(\logo_left[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2636_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0038_),
    .Q(\logo_left[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2637_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0039_),
    .Q(\logo_left[8] ));
 sky130_fd_sc_hd__dfxtp_2 _2638_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0040_),
    .Q(\logo_left[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2639_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0041_),
    .Q(\logo_top[0] ));
 sky130_fd_sc_hd__dfxtp_4 _2640_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0042_),
    .Q(\logo_top[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2641_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0043_),
    .Q(\logo_top[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2642_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0044_),
    .Q(\logo_top[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2643_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0045_),
    .Q(\logo_top[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2644_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0046_),
    .Q(\logo_top[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2645_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0047_),
    .Q(\logo_top[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2646_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0048_),
    .Q(\logo_top[7] ));
 sky130_fd_sc_hd__dfxtp_2 _2647_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0049_),
    .Q(\logo_top[8] ));
 sky130_fd_sc_hd__dfxtp_2 _2648_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0050_),
    .Q(\logo_top[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2649_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0051_),
    .Q(dir_x));
 sky130_fd_sc_hd__dfxtp_1 _2650_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0052_),
    .Q(dir_y));
 sky130_fd_sc_hd__dfxtp_1 _2651_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0053_),
    .Q(manual_mode));
 sky130_fd_sc_hd__dfxtp_1 _2652_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0054_),
    .Q(\color_index[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2653_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0055_),
    .Q(\color_index[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2654_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0056_),
    .Q(\color_index[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2655_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0057_),
    .Q(\prev_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2656_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0058_),
    .Q(\prev_y[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2657_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0059_),
    .Q(\prev_y[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2658_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0060_),
    .Q(\prev_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2659_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0061_),
    .Q(\prev_y[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2660_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0062_),
    .Q(\prev_y[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2661_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0063_),
    .Q(\prev_y[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2662_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0064_),
    .Q(\prev_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2663_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0065_),
    .Q(\prev_y[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2664_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0066_),
    .Q(\prev_y[9] ));
 sky130_fd_sc_hd__dfxtp_2 _2665_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0067_),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__dfxtp_2 _2666_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0068_),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__dfxtp_2 _2667_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0069_),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__dfxtp_2 _2668_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0070_),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__dfxtp_1 _2669_ (.CLK(clknet_3_4__leaf_clk),
    .D(net154),
    .Q(\gamepad.driver.pmod_clk_prev ));
 sky130_fd_sc_hd__dfxtp_1 _2670_ (.CLK(clknet_3_4__leaf_clk),
    .D(net155),
    .Q(\gamepad.driver.pmod_latch_prev ));
 sky130_fd_sc_hd__dfxtp_1 _2671_ (.CLK(clknet_3_4__leaf_clk),
    .D(net172),
    .Q(\gamepad.driver.shift_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2672_ (.CLK(clknet_3_4__leaf_clk),
    .D(net192),
    .Q(\gamepad.driver.shift_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2673_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0073_),
    .Q(\gamepad.driver.shift_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2674_ (.CLK(clknet_3_7__leaf_clk),
    .D(net179),
    .Q(\gamepad.driver.shift_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2675_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0075_),
    .Q(\gamepad.driver.shift_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2676_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0076_),
    .Q(\gamepad.driver.shift_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2677_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0077_),
    .Q(\gamepad.driver.shift_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2678_ (.CLK(clknet_3_6__leaf_clk),
    .D(net185),
    .Q(\gamepad.driver.shift_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2679_ (.CLK(clknet_3_7__leaf_clk),
    .D(net181),
    .Q(\gamepad.driver.shift_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2680_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0080_),
    .Q(\gamepad.driver.shift_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2681_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0081_),
    .Q(\gamepad.driver.shift_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2682_ (.CLK(clknet_3_7__leaf_clk),
    .D(net177),
    .Q(\gamepad.driver.shift_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2683_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0083_),
    .Q(\gamepad.driver.pmod_data_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2684_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0084_),
    .Q(\gamepad.driver.pmod_data_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2685_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0085_),
    .Q(\gamepad.driver.pmod_clk_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2686_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0086_),
    .Q(\gamepad.driver.pmod_clk_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2687_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0087_),
    .Q(\gamepad.driver.pmod_latch_sync[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2688_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0088_),
    .Q(\gamepad.driver.pmod_latch_sync[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2689_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0004_),
    .Q(hsync));
 sky130_fd_sc_hd__dfxtp_2 _2690_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0089_),
    .Q(\pix_y[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2691_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0090_),
    .Q(\pix_y[1] ));
 sky130_fd_sc_hd__dfxtp_2 _2692_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0091_),
    .Q(\pix_y[2] ));
 sky130_fd_sc_hd__dfxtp_2 _2693_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0092_),
    .Q(\pix_y[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2694_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0093_),
    .Q(\pix_y[4] ));
 sky130_fd_sc_hd__dfxtp_2 _2695_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0094_),
    .Q(\pix_y[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2696_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0095_),
    .Q(\pix_y[6] ));
 sky130_fd_sc_hd__dfxtp_2 _2697_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0096_),
    .Q(\pix_y[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2698_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0097_),
    .Q(\pix_y[8] ));
 sky130_fd_sc_hd__dfxtp_2 _2699_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0098_),
    .Q(\pix_y[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2700_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0005_),
    .Q(\vga_sync_gen.vsync ));
 sky130_fd_sc_hd__dfxtp_1 _2701_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0099_),
    .Q(\palette_inst.rrggbb[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2702_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0000_),
    .Q(\palette_inst.rrggbb[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2703_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0001_),
    .Q(\palette_inst.rrggbb[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2704_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0002_),
    .Q(\palette_inst.rrggbb[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2705_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0003_),
    .Q(\palette_inst.rrggbb[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2706_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0100_),
    .Q(\palette_inst.rrggbb[4] ));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_139 (.LO(net139));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_140 (.LO(net140));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_141 (.LO(net141));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_142 (.LO(net142));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_143 (.LO(net143));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_144 (.LO(net144));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_145 (.LO(net145));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_146 (.LO(net146));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_147 (.LO(net147));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_148 (.LO(net148));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_149 (.LO(net149));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_150 (.LO(net150));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_151 (.LO(net151));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_152 (.LO(net152));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_153 (.LO(net153));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__buf_2 _2723_ (.A(\vga_sync_gen.vsync ),
    .X(uo_out[3]));
 sky130_fd_sc_hd__buf_2 _2724_ (.A(hsync),
    .X(uo_out[7]));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_617 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 wire7 (.A(_1064_),
    .X(net7));
 sky130_fd_sc_hd__buf_4 fanout8 (.A(_0624_),
    .X(net8));
 sky130_fd_sc_hd__buf_2 fanout9 (.A(_0383_),
    .X(net9));
 sky130_fd_sc_hd__buf_2 fanout10 (.A(_0258_),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout11 (.A(_0258_),
    .X(net11));
 sky130_fd_sc_hd__buf_2 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 fanout14 (.A(_0760_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(_0759_),
    .X(net16));
 sky130_fd_sc_hd__buf_2 fanout17 (.A(_0726_),
    .X(net17));
 sky130_fd_sc_hd__buf_2 fanout18 (.A(_0712_),
    .X(net18));
 sky130_fd_sc_hd__buf_2 fanout19 (.A(net20),
    .X(net19));
 sky130_fd_sc_hd__buf_4 fanout20 (.A(_0682_),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout21 (.A(_0667_),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(_0663_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout23 (.A(net25),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(_0658_),
    .X(net25));
 sky130_fd_sc_hd__buf_2 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(net29),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(_0657_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(_0750_),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_4 fanout31 (.A(_0741_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_4 fanout33 (.A(_0738_),
    .X(net33));
 sky130_fd_sc_hd__buf_4 fanout34 (.A(_0720_),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_4 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(_0719_),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(_0706_),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 fanout40 (.A(_0705_),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(_0705_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(_0688_),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net49),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(net49),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net49),
    .X(net46));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout47 (.A(net49),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_2 fanout49 (.A(_0661_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net54),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(net54),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(_0660_),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(_0656_),
    .X(net55));
 sky130_fd_sc_hd__buf_2 fanout56 (.A(net57),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 fanout57 (.A(_0656_),
    .X(net57));
 sky130_fd_sc_hd__buf_2 fanout58 (.A(_0655_),
    .X(net58));
 sky130_fd_sc_hd__buf_2 fanout59 (.A(_0655_),
    .X(net59));
 sky130_fd_sc_hd__buf_2 fanout60 (.A(_0654_),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(_0654_),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_4 fanout63 (.A(net65),
    .X(net63));
 sky130_fd_sc_hd__buf_2 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 fanout65 (.A(_0653_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(_0631_),
    .X(net66));
 sky130_fd_sc_hd__buf_2 fanout67 (.A(_0631_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(_0833_),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(_0731_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(net72),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__buf_2 fanout72 (.A(_0730_),
    .X(net72));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(_0687_),
    .X(net73));
 sky130_fd_sc_hd__buf_2 fanout74 (.A(_0686_),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(_0676_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_8 fanout76 (.A(_0675_),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(net78),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(_0665_),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_8 fanout79 (.A(_0664_),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(_0664_),
    .X(net80));
 sky130_fd_sc_hd__buf_4 fanout81 (.A(_0627_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 fanout82 (.A(_0627_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(_0627_),
    .X(net83));
 sky130_fd_sc_hd__buf_2 fanout84 (.A(_0627_),
    .X(net84));
 sky130_fd_sc_hd__buf_4 fanout85 (.A(_0626_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 fanout86 (.A(_0626_),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_4 fanout87 (.A(net89),
    .X(net87));
 sky130_fd_sc_hd__buf_2 fanout88 (.A(net89),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(_0626_),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(_0685_),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(_0685_),
    .X(net91));
 sky130_fd_sc_hd__buf_2 fanout92 (.A(_0685_),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(_0685_),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(_0684_),
    .X(net94));
 sky130_fd_sc_hd__buf_2 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(_0684_),
    .X(net97));
 sky130_fd_sc_hd__buf_4 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(_0629_),
    .X(net99));
 sky130_fd_sc_hd__buf_4 fanout100 (.A(net102),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(net102),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(_0628_),
    .X(net102));
 sky130_fd_sc_hd__buf_2 fanout103 (.A(_0491_),
    .X(net103));
 sky130_fd_sc_hd__buf_2 fanout104 (.A(_0244_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(net108),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(net108),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(net108),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(_0633_),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(_0632_),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 fanout112 (.A(_0632_),
    .X(net112));
 sky130_fd_sc_hd__buf_2 fanout113 (.A(_0490_),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(_0243_),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(_0518_),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(_0517_),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(_0516_),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(\pix_y[8] ),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_4 fanout119 (.A(\pix_y[1] ),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(manual_mode),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(manual_mode),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(manual_mode),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(manual_mode),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(dir_y),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_4 fanout125 (.A(\logo_top[7] ),
    .X(net125));
 sky130_fd_sc_hd__buf_2 fanout126 (.A(\logo_top[6] ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(\logo_top[5] ),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_2 fanout128 (.A(\logo_top[4] ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(\logo_top[3] ),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(\logo_left[4] ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 fanout131 (.A(\logo_left[3] ),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net137),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net137),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout134 (.A(net137),
    .X(net134));
 sky130_fd_sc_hd__buf_2 fanout135 (.A(net137),
    .X(net135));
 sky130_fd_sc_hd__buf_1 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net1),
    .X(net137));
 sky130_fd_sc_hd__conb_1 tt_um_zerotoasic_logo_screensaver_138 (.LO(net138));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload2 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\gamepad.driver.pmod_clk_sync[1] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\gamepad.driver.pmod_latch_sync[1] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\gamepad.driver.pmod_latch_sync[0] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\gamepad.driver.pmod_data_sync[0] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\gamepad.driver.pmod_clk_sync[0] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\gamepad.decoder.data_reg[11] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0019_),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\gamepad.decoder.data_reg[2] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0010_),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\gamepad.decoder.data_reg[0] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_0008_),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\gamepad.decoder.data_reg[9] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0017_),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\gamepad.decoder.data_reg[1] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_0009_),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\gamepad.decoder.data_reg[10] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0018_),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\gamepad.driver.pmod_data_sync[1] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0071_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\gamepad.decoder.data_reg[3] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_0011_),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\palette_inst.rrggbb[5] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\gamepad.driver.shift_reg[11] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0082_),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\gamepad.driver.shift_reg[3] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0074_),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\gamepad.driver.shift_reg[8] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0079_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\palette_inst.rrggbb[3] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\gamepad.driver.shift_reg[4] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\gamepad.driver.shift_reg[7] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0078_),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\gamepad.driver.shift_reg[5] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\gamepad.decoder.data_reg[8] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\gamepad.driver.shift_reg[6] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\gamepad.driver.shift_reg[9] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\gamepad.driver.shift_reg[10] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\gamepad.driver.shift_reg[1] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0072_),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\prev_y[5] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\gamepad.decoder.data_reg[5] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\prev_y[9] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\prev_y[4] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\gamepad.decoder.data_reg[4] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\gamepad.decoder.data_reg[6] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\gamepad.driver.shift_reg[2] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\prev_y[6] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\prev_y[8] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\prev_y[0] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\prev_y[3] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\prev_y[7] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\prev_y[2] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\color_index[1] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\gamepad.decoder.data_reg[7] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\pix_x[2] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\prev_y[1] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\logo_left[0] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\pix_x[9] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\pix_x[0] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\pix_x[5] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\pix_y[3] ),
    .X(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__D (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1328__X (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__D (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1325__X (.DIODE(_0005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A3 (.DIODE(_0157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__X (.DIODE(_0157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2382__B1 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__A (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__B1 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2306__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__A2 (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__Y (.DIODE(_0280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__C1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__C1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2417__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__C1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__C1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__C1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__C1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2271__A (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__A (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__Y (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2181__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__B2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__B2 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__Y (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2304__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2303__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__S (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__B (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1343__X (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__B (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__B (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__X (.DIODE(_0586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_A (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__A1 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1421__X (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__B1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__A1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__C1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1935__C1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__C1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A1 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__Y (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__X (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1424__Y (.DIODE(_0627_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__B1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__Y (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__C1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A1_N (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1932__A (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A1_N (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__A1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__B1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__B2 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__B1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__B1 (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__Y (.DIODE(_0630_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__X (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__A1 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1451__Y (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__B (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__A2 (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1453__X (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__A_N (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__B1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__X (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__C1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__D1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__X (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__A2 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1663__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1510__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__X (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__S (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A1 (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__X (.DIODE(_0684_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__Y (.DIODE(_0685_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__A2 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__A1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__B2 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__Y (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A3 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__X (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__B2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__B2 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1709__A1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__A2_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__X (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__B2 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A3 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__C_N (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__B1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__B1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__C1 (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__Y (.DIODE(_0699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A1_N (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__C1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__X (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A1 (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__X (.DIODE(_0705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__A (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__B2 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__A (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__Y (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__A (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__A (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__A1 (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1508__Y (.DIODE(_0711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__A (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__C (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1576__A2 (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__A (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__Y (.DIODE(_0714_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__C1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__A1 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__B2 (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__Y (.DIODE(_0720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__B2 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__B1 (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__A (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__Y (.DIODE(_0722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__B2 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__B (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A_N (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A1 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__A2 (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__C (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__B (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__B (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__X (.DIODE(_0728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__A (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__X (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__C1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A1 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__A (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__A2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__A2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__A2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__A2 (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__B (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__X (.DIODE(_0732_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A1 (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__Y (.DIODE(_0738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__B2 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__B1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__B (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__A1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__B1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__B1 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__Y (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__B2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__C (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__B1 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__Y (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__B (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__B2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__B1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__A2 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__X (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__B2 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__C1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__C1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1592__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__B (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__Y (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__A2 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1552__A2 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__X (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__A1 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__A2 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__A2 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__C (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__A2 (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__B (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__C (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__Y (.DIODE(_0762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__B (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A2 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__C (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__Y (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1795__A1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__B (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__B (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__A1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__Y (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__B1 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__A1 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2096__B (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__B (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__A3 (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__B (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__B (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__Y (.DIODE(_0778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__A (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__A2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__A2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__A1 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__A2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A2 (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1712__B (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__A2_N (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__B (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__Y (.DIODE(_0790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__B1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__B1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__A2 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1843__B1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__A2 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__Y (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__B (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__B1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__A1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1845__B (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A2 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__C (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__B1 (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1596__B (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__Y (.DIODE(_0798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__B (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__A2 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A2 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__Y (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A2 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__A2 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__B1 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A3 (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__X (.DIODE(_0828_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__Y (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A2 (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A2 (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A3 (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__B (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1831__A (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__Y (.DIODE(_0834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2135__A (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__Y (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__A2 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1806__A1 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__A2 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__A2 (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__X (.DIODE(_0840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__B1 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__B1 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__B1 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__B1 (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__A (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__Y (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1906__A2 (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A1 (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__A (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__A1 (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__X (.DIODE(_0847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__C1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__B1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__A (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__B1 (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__B (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__B (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__Y (.DIODE(_0850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__A (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__B (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__B1 (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__B (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__Y (.DIODE(_0851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__C1 (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__Y (.DIODE(_0852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__B1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__B1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__B (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__B1 (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__Y (.DIODE(_0853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__B2 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__A2 (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__A (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__Y (.DIODE(_0864_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__A1 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__A2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__B2 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__C1 (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__Y (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1915__A2 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1823__A3 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__A1 (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__X (.DIODE(_0873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__B1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__A2 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__B1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__A1 (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__Y (.DIODE(_0878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__A1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__B2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__A2 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__B1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__B1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__B1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__B1 (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__Y (.DIODE(_0879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__B1 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__B (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__B (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A2 (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1680__X (.DIODE(_0883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__A1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__B1 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__A3 (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__X (.DIODE(_0898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__C (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__B (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__B2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__A2 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__A0 (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__B (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__Y (.DIODE(_0901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__B1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A3 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__B2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A3 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__B (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__A3 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__X (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__B2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__Y (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__A2 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__B1 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2102__A2 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__A2 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A3 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A2 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A2 (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__X (.DIODE(_0945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A1 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2019__A3 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A2 (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__C (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__Y (.DIODE(_0947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__A (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__A2 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A2 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__B2 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A2 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__B1 (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__Y (.DIODE(_0950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__A2 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2160__B1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__B1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__B2 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__B2 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__A1 (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__Y (.DIODE(_0951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A2 (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__Y (.DIODE(_0959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__A2 (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A2_N (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2041__B (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A_N (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__B1 (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__Y (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__B1 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__B1 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__A1 (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__Y (.DIODE(_0971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__B2 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__A1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A2 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1803__B1 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1800__A2 (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__Y (.DIODE(_0972_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__B (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__A (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__B1 (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__A2 (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__Y (.DIODE(_0976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__C1 (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__X (.DIODE(_0991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__B2 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2082__A (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__D1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__Y (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__B1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__B1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__B1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__C1 (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__Y (.DIODE(_1037_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__A2 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__B (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__A1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__C (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__A2 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__B1 (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__Y (.DIODE(_1076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A3 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A4 (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__X (.DIODE(_1079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__B1 (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__B1 (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__Y (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__A2 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__C (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__A1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A2 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__B1 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__X (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__A2 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__X (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__S (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__B2 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1916__A2 (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__Y (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__B2 (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__X (.DIODE(_1247_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__Q (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__A (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A1 (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A1 (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A1 (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__B (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__A2 (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__B (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1331__A (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__A (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__A (.DIODE(\pix_y[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__Q (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A1 (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B1 (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A1 (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__B (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__B (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1340__C (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__A (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B (.DIODE(\pix_y[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__Q (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A1 (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__A_N (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__B (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A1 (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__B (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__2179__B (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__D (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__A (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__B_N (.DIODE(\pix_y[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(ui_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(ui_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(ui_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(ui_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(ui_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_X (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1722__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__C1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__C1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1657__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__C1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_X (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__B (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A0 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_X (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__C1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1598__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__C1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_X (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__C1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1787__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__C1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_X (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__C1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__C1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1801__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__C1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__C1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1721__C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__C1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1788__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_X (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__C1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__C1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_X (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1807__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1851__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__C1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_X (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1662__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1848__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1588__A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__A1_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__S0 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_X (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__2124__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__2061__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2075__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_X (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1850__B1_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1580__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1914__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__C1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A2_N (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_X (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__A1_N (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__C1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__A3 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2139__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__A1_N (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_X (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1796__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2013__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1606__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__2033__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1790__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1907__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__C1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1638__C1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_X (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__C1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2157__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__C1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A1_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__C1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_X (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__C1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__2079__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1708__C1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__1934__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_X (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__C1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__C1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_X (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__D1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2074__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__C1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__1624__C1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__C1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__C1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__C1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_X (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__D1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1799__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__C1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__B (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__C1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__C1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__1852__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_X (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__C1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1703__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__C (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__C1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1626__A0 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A3 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1467__C (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1550__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1586__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1582__A1_N (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_X (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_X (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__S (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__B1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1716__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__C (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_X (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__S (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1636__A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_X (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_X (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__B (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1455__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1717__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_X (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__C1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_X (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__1454__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__2186__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1710__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__C1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__C1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_X (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__2084__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__C1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__B (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_X (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1843__A2_N (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__B (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1608__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__2159__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_X (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_X (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2168__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1853__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1572__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1842__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__2158__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_X (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__B (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1590__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_X (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2222__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__D (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__B (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1566__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__C1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__D (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1568__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__B (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_X (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__A3 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__B (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__C1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__C (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1562__C1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__D (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_X (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1680__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1464__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__C1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__C (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__1570__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_X (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1797__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__1713__C1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__C1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__D1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_X (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1714__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__C1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1821__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__D1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__1827__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__1805__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__1804__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__D1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_X (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1578__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1809__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__B2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1798__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__1794__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__C1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_X (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__C (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_X (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__D1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__B (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1802__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_X (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1793__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__B (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__2144__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_X (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__1546__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__S1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_X (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__B (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1820__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__2146__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_X (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__1427__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1634__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__2076__C1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__B (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_X (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_X (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__C1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__B (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__1720__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_X (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__C1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2156__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1639__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1594__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__1709__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__2072__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1789__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_X (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__C1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__C1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1893__C1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1574__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1844__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1622__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__B (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_X (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2312__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2328__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2384__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2388__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_X (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2326__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2473__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__2436__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__C (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2180__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__D (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1342__B (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2489__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_X (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2354__S (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2349__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__A_N (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_X (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2263__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1319__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2471__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2461__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__C1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_X (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1387__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__C1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2305__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_X (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__C1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__CLK (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_X (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1065_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0145_));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_299 ();
 assign uio_oe[0] = net138;
 assign uio_oe[1] = net139;
 assign uio_oe[2] = net140;
 assign uio_oe[3] = net141;
 assign uio_oe[4] = net142;
 assign uio_oe[5] = net143;
 assign uio_oe[6] = net144;
 assign uio_oe[7] = net145;
 assign uio_out[0] = net146;
 assign uio_out[1] = net147;
 assign uio_out[2] = net148;
 assign uio_out[3] = net149;
 assign uio_out[4] = net150;
 assign uio_out[5] = net151;
 assign uio_out[6] = net152;
 assign uio_out[7] = net153;
endmodule
